*SPICE netlist created from verilog structural netlist module atbs_core_floating_window_board by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

.subckt atbs_core_floating_window_board VPWR VGND adaptive_mode_i clock_i comp_lower_i comp_upper_i control_mode_i
+ dac_lower_o[0] dac_lower_o[1] dac_lower_o[2] dac_lower_o[3] dac_lower_o[4] dac_lower_o[5] dac_lower_o[6] dac_lower_o[7]
+ dac_upper_o[0] dac_upper_o[1] dac_upper_o[2] dac_upper_o[3] dac_upper_o[4] dac_upper_o[5] dac_upper_o[6] dac_upper_o[7]
+ enable_i idle_led_o overflow_led_o reset_n_i select_tbs_delta_steps_i signal_select_in_i trigger_start_mode_i trigger_start_sampling_i
+ uart_rx_i uart_tx_o underflow_led_o 

X_06941_ \atbs_core_0.uart_0.uart_rx_0.n2848_o\ VPWR VGND _00748_ sg13g2_buf_1
X_06942_ _00748_ VPWR VGND _00749_ sg13g2_inv_1
X_06943_ \atbs_core_0.baudrate_adj_uart[2]\ VPWR VGND _00750_ sg13g2_buf_1
X_06944_ _00750_ VPWR VGND _00751_ sg13g2_inv_1
X_06945_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[2]\ VPWR VGND _00752_ sg13g2_buf_1
X_06946_ \atbs_core_0.baudrate_adj_uart[5]\ VPWR VGND _00753_ sg13g2_buf_1
X_06947_ _00753_ VPWR VGND _00754_ sg13g2_buf_1
X_06948_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[5]\ VPWR VGND _00755_ sg13g2_buf_1
X_06949_ _00754_ _00755_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ VPWR VGND _00756_ sg13g2_nand3_1
X_06950_ _00753_ _00755_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ VPWR VGND _00757_ sg13g2_or3_1
X_06951_ \atbs_core_0.baudrate_adj_uart[6]\ VPWR VGND _00758_ sg13g2_buf_1
X_06952_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[6]\ VPWR VGND _00759_ sg13g2_buf_1
X_06953_ _00758_ _00759_ VPWR VGND _00760_ sg13g2_xor2_1
X_06954_ _00751_ _00752_ _00756_ _00757_ _00760_ VPWR 
+ VGND
+ _00761_ sg13g2_a221oi_1
X_06955_ \atbs_core_0.baudrate_adj_uart[4]\ VPWR VGND _00762_ sg13g2_buf_1
X_06956_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[4]\ VPWR VGND _00763_ sg13g2_buf_1
X_06957_ _00762_ _00763_ VPWR VGND _00764_ sg13g2_nand2b_1
X_06958_ _00763_ _00762_ VPWR VGND _00765_ sg13g2_nand2b_1
X_06959_ _00752_ VPWR VGND _00766_ sg13g2_inv_1
X_06960_ \atbs_core_0.baudrate_adj_uart[1]\ VPWR VGND _00767_ sg13g2_buf_1
X_06961_ _00767_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ VPWR VGND _00768_ sg13g2_xor2_1
X_06962_ _00750_ _00766_ _00768_ VPWR VGND _00769_ sg13g2_a21oi_1
X_06963_ _00764_ _00765_ _00769_ VPWR VGND _00770_ sg13g2_and3_1
X_06964_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[1]\ VPWR VGND _00771_ sg13g2_buf_1
X_06965_ _00767_ _00771_ VPWR VGND _00772_ sg13g2_xor2_1
X_06966_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[0]\ VPWR VGND _00773_ sg13g2_buf_1
X_06967_ \atbs_core_0.baudrate_adj_uart[0]\ VPWR VGND _00774_ sg13g2_buf_1
X_06968_ _00773_ _00774_ VPWR VGND _00775_ sg13g2_xor2_1
X_06969_ \atbs_core_0.baudrate_adj_uart[7]\ VPWR VGND _00776_ sg13g2_buf_1
X_06970_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ VPWR VGND _00777_ sg13g2_buf_1
X_06971_ _00777_ VPWR VGND _00778_ sg13g2_inv_1
X_06972_ _00776_ _00778_ VPWR VGND _00779_ sg13g2_nor2_1
X_06973_ _00776_ VPWR VGND _00780_ sg13g2_inv_1
X_06974_ _00780_ _00777_ VPWR VGND _00781_ sg13g2_nor2_1
X_06975_ _00772_ _00775_ _00779_ _00781_ VPWR VGND 
+ _00782_
+ sg13g2_nor4_1
X_06976_ _00761_ _00770_ _00782_ VPWR VGND _00783_ sg13g2_nand3_1
X_06977_ _00783_ VPWR VGND _00784_ sg13g2_buf_1
X_06978_ \atbs_core_0.uart_0.uart_rx_0.n2891_o\ VPWR VGND _00785_ sg13g2_buf_1
X_06979_ \atbs_core_0.uart_0.uart_rx_0.n2889_o\ VPWR VGND _00786_ sg13g2_buf_1
X_06980_ \atbs_core_0.uart_0.uart_rx_0.n2897_o\ VPWR VGND _00787_ sg13g2_buf_1
X_06981_ _00785_ _00786_ _00787_ VPWR VGND _00788_ sg13g2_nand3_1
X_06982_ \atbs_core_0.uart_0.uart_rx_0.n2819_o\ VPWR VGND _00789_ sg13g2_buf_1
X_06983_ _00784_ _00788_ _00789_ VPWR VGND _00790_ sg13g2_o21ai_1
X_06984_ _00749_ _00784_ _00790_ VPWR VGND _00000_ sg13g2_o21ai_1
X_06985_ \atbs_core_0.uart_0.uart_tx_0.n2735_o\ VPWR VGND _00791_ sg13g2_buf_1
X_06986_ _00791_ VPWR VGND _00792_ sg13g2_inv_1
X_06987_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[7]\ VPWR VGND _00793_ sg13g2_buf_1
X_06988_ _00776_ _00793_ VPWR VGND _00794_ sg13g2_xnor2_1
X_06989_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[4]\ VPWR VGND _00795_ sg13g2_buf_1
X_06990_ _00762_ _00795_ VPWR VGND _00796_ sg13g2_xnor2_1
X_06991_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[5]\ VPWR VGND _00797_ sg13g2_buf_1
X_06992_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[8]\ VPWR VGND _00798_ sg13g2_buf_1
X_06993_ _00754_ _00797_ _00798_ VPWR VGND _00799_ sg13g2_nand3_1
X_06994_ _00753_ _00797_ _00798_ VPWR VGND _00800_ sg13g2_or3_1
X_06995_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[1]\ VPWR VGND _00801_ sg13g2_buf_1
X_06996_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[3]\ VPWR VGND _00802_ sg13g2_buf_1
X_06997_ _00767_ _00801_ _00802_ VPWR VGND _00803_ sg13g2_or3_1
X_06998_ _00767_ _00801_ _00802_ VPWR VGND _00804_ sg13g2_nand3_1
X_06999_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[2]\ VPWR VGND _00805_ sg13g2_buf_1
X_07000_ _00751_ _00805_ VPWR VGND _00806_ sg13g2_nand2_1
X_07001_ _00805_ _00750_ VPWR VGND _00807_ sg13g2_nand2b_1
X_07002_ _00758_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ VPWR VGND _00808_ sg13g2_xnor2_1
X_07003_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[0]\ VPWR VGND _00809_ sg13g2_buf_1
X_07004_ _00774_ _00809_ VPWR VGND _00810_ sg13g2_xnor2_1
X_07005_ _00806_ _00807_ _00808_ _00810_ VPWR VGND 
+ _00811_
+ sg13g2_nand4_1
X_07006_ _00799_ _00800_ _00803_ _00804_ _00811_ VPWR 
+ VGND
+ _00812_ sg13g2_a221oi_1
X_07007_ _00794_ _00796_ _00812_ VPWR VGND _00813_ sg13g2_nand3_1
X_07008_ _00813_ VPWR VGND _00814_ sg13g2_buf_1
X_07009_ _00814_ VPWR VGND _00815_ sg13g2_buf_1
X_07010_ \atbs_core_0.uart_0.uart_tx_0.n2730_o\ VPWR VGND _00816_ sg13g2_buf_1
X_07011_ \atbs_core_0.uart_0.uart_tx_0.n2758_o\ VPWR VGND _00817_ sg13g2_inv_1
X_07012_ \atbs_core_0.uart_0.uart_tx_0.n2721_o\ VPWR VGND _00818_ sg13g2_inv_1
X_07013_ \atbs_core_0.memory2uart_0.n2040_q\ VPWR VGND _00819_ sg13g2_inv_1
X_07014_ _00817_ _00818_ _00819_ VPWR VGND _00820_ sg13g2_a21oi_1
X_07015_ _00816_ _00815_ _00820_ VPWR VGND _00821_ sg13g2_nor3_1
X_07016_ _00792_ _00815_ _00821_ VPWR VGND _00003_ sg13g2_a21oi_1
X_07017_ _00028_ VPWR VGND _00822_ sg13g2_inv_1
X_07018_ \atbs_core_0.dac_control_0.n1586_q\ VPWR VGND _00823_ sg13g2_buf_1
X_07019_ _00823_ VPWR VGND _00824_ sg13g2_inv_1
X_07020_ \atbs_core_0.main_counter_value[5]\ VPWR VGND _00825_ sg13g2_buf_1
X_07021_ \atbs_core_0.main_counter_value[2]\ _00825_ \atbs_core_0.main_counter_value[7]\ \atbs_core_0.main_counter_value[6]\ VPWR VGND 
+ _00826_
+ sg13g2_nor4_1
X_07022_ \atbs_core_0.main_counter_value[9]\ VPWR VGND _00827_ sg13g2_buf_1
X_07023_ \atbs_core_0.main_counter_value[8]\ VPWR VGND _00828_ sg13g2_buf_1
X_07024_ \atbs_core_0.main_counter_value[17]\ VPWR VGND _00829_ sg13g2_buf_1
X_07025_ \atbs_core_0.main_counter_value[16]\ VPWR VGND _00830_ sg13g2_buf_1
X_07026_ \atbs_core_0.main_counter_value[15]\ \atbs_core_0.main_counter_value[14]\ _00829_ _00830_ VPWR VGND 
+ _00831_
+ sg13g2_or4_1
X_07027_ _00827_ _00828_ \atbs_core_0.main_counter_value[11]\ _00831_ VPWR VGND 
+ _00832_
+ sg13g2_nor4_1
X_07028_ \atbs_core_0.main_counter_value[18]\ VPWR VGND _00833_ sg13g2_buf_1
X_07029_ _00833_ \atbs_core_0.main_counter_value[19]\ VPWR VGND _00834_ sg13g2_nor2_1
X_07030_ \atbs_core_0.main_counter_value[0]\ VPWR VGND _00835_ sg13g2_buf_1
X_07031_ \atbs_core_0.main_counter_value[10]\ VPWR VGND _00836_ sg13g2_buf_1
X_07032_ \atbs_core_0.main_counter_value[13]\ VPWR VGND _00837_ sg13g2_buf_1
X_07033_ \atbs_core_0.main_counter_value[12]\ VPWR VGND _00838_ sg13g2_buf_1
X_07034_ _00835_ _00836_ _00837_ _00838_ VPWR VGND 
+ _00839_
+ sg13g2_nor4_1
X_07035_ _00826_ _00832_ _00834_ _00839_ VPWR VGND 
+ _00840_
+ sg13g2_and4_1
X_07036_ _00840_ VPWR VGND _00841_ sg13g2_buf_1
X_07037_ \atbs_core_0.n1074_q[2]\ VPWR VGND _00842_ sg13g2_buf_1
X_07038_ \atbs_core_0.n1074_q[0]\ VPWR VGND _00843_ sg13g2_buf_1
X_07039_ _00843_ VPWR VGND _00844_ sg13g2_inv_1
X_07040_ _00844_ _00027_ VPWR VGND _00845_ sg13g2_nand2_1
X_07041_ \atbs_core_0.main_counter_value[1]\ VPWR VGND _00846_ sg13g2_buf_1
X_07042_ \atbs_core_0.main_counter_value[3]\ VPWR VGND _00847_ sg13g2_inv_1
X_07043_ \atbs_core_0.main_counter_value[4]\ VPWR VGND _00848_ sg13g2_buf_1
X_07044_ \atbs_core_0.n1074_q[1]\ VPWR VGND _00849_ sg13g2_buf_1
X_07045_ _00846_ _00847_ _00848_ _00849_ VPWR VGND 
+ _00850_
+ sg13g2_nand4_1
X_07046_ _00842_ _00845_ _00850_ VPWR VGND _00851_ sg13g2_nor3_1
X_07047_ _00841_ _00851_ VPWR VGND _00852_ sg13g2_nand2_1
X_07048_ \atbs_core_0.control_mode_debounced\ VPWR VGND _00853_ sg13g2_buf_16
X_07049_ _00853_ _00008_ VPWR VGND _00854_ sg13g2_nor2b_1
X_07050_ _00009_ _00853_ _00854_ VPWR VGND _00855_ sg13g2_a21oi_2
X_07051_ _00855_ VPWR VGND _00856_ sg13g2_buf_1
X_07052_ _00856_ VPWR VGND _00857_ sg13g2_buf_1
X_07053_ _00857_ VPWR VGND _00858_ sg13g2_buf_1
X_07054_ _00024_ VPWR VGND _00859_ sg13g2_buf_1
X_07055_ \atbs_core_0.adaptive_ctrl_0.adapt_on_overflow\ VPWR VGND _00860_ sg13g2_buf_2
X_07056_ _00860_ VPWR VGND _00861_ sg13g2_inv_1
X_07057_ _00861_ VPWR VGND _00862_ sg13g2_buf_1
X_07058_ _00025_ VPWR VGND _00863_ sg13g2_inv_1
X_07059_ \atbs_core_0.spike_detector_0.lock_detection\ \atbs_core_0.detection_en\ VPWR VGND _00864_ sg13g2_nand2b_1
X_07060_ _00008_ _00009_ _00853_ VPWR VGND _00865_ sg13g2_mux2_1
X_07061_ _00865_ VPWR VGND _00866_ sg13g2_buf_4
X_07062_ \atbs_core_0.n1054_q\ _00866_ VPWR VGND _00867_ sg13g2_nor2b_2
X_07063_ \atbs_core_0.adaptive_ctrl_0.n1373_o[5]\ VPWR VGND _00868_ sg13g2_buf_1
X_07064_ \atbs_core_0.adaptive_ctrl_0.n1373_o[4]\ VPWR VGND _00869_ sg13g2_buf_2
X_07065_ _00868_ _00869_ VPWR VGND _00870_ sg13g2_or2_1
X_07066_ \atbs_core_0.adaptive_ctrl_0.n1373_o[1]\ VPWR VGND _00871_ sg13g2_buf_4
X_07067_ \atbs_core_0.adaptive_ctrl_0.n1373_o[0]\ VPWR VGND _00872_ sg13g2_buf_2
X_07068_ \atbs_core_0.adaptive_ctrl_0.n1373_o[6]\ VPWR VGND _00873_ sg13g2_buf_2
X_07069_ \atbs_core_0.adaptive_ctrl_0.n1449_q[8]\ VPWR VGND _00874_ sg13g2_buf_2
X_07070_ _00871_ _00872_ _00873_ _00874_ VPWR VGND 
+ _00875_
+ sg13g2_or4_1
X_07071_ \atbs_core_0.adaptive_ctrl_0.n1373_o[3]\ VPWR VGND _00876_ sg13g2_buf_2
X_07072_ \atbs_core_0.adaptive_ctrl_0.n1373_o[2]\ VPWR VGND _00877_ sg13g2_buf_1
X_07073_ \atbs_core_0.adaptive_ctrl_0.n1373_o[7]\ VPWR VGND _00878_ sg13g2_buf_2
X_07074_ _00876_ _00877_ _00878_ VPWR VGND _00879_ sg13g2_or3_1
X_07075_ _00866_ _00870_ _00875_ _00879_ VPWR VGND 
+ _00880_
+ sg13g2_nor4_2
X_07076_ \atbs_core_0.comp_lower_sync\ _00864_ _00867_ _00880_ VPWR VGND 
+ _00881_
+ sg13g2_or4_1
X_07077_ _00881_ VPWR VGND _00882_ sg13g2_buf_8
X_07078_ _00866_ VPWR VGND _00883_ sg13g2_buf_16
X_07079_ \atbs_core_0.adaptive_ctrl_0.n1368_o[7]\ VPWR VGND _00884_ sg13g2_buf_1
X_07080_ \atbs_core_0.adaptive_ctrl_0.n1448_q[8]\ VPWR VGND _00885_ sg13g2_buf_1
X_07081_ _00884_ _00885_ VPWR VGND _00886_ sg13g2_or2_1
X_07082_ \atbs_core_0.adaptive_ctrl_0.n1368_o[1]\ VPWR VGND _00887_ sg13g2_buf_1
X_07083_ \atbs_core_0.adaptive_ctrl_0.n1368_o[5]\ VPWR VGND _00888_ sg13g2_buf_1
X_07084_ \atbs_core_0.adaptive_ctrl_0.n1368_o[4]\ VPWR VGND _00889_ sg13g2_buf_1
X_07085_ \atbs_core_0.adaptive_ctrl_0.n1368_o[6]\ VPWR VGND _00890_ sg13g2_buf_2
X_07086_ _00887_ _00888_ _00889_ _00890_ VPWR VGND 
+ _00891_
+ sg13g2_or4_1
X_07087_ \atbs_core_0.adaptive_ctrl_0.n1368_o[0]\ VPWR VGND _00892_ sg13g2_buf_2
X_07088_ \atbs_core_0.adaptive_ctrl_0.n1368_o[3]\ VPWR VGND _00893_ sg13g2_buf_2
X_07089_ \atbs_core_0.adaptive_ctrl_0.n1368_o[2]\ VPWR VGND _00894_ sg13g2_buf_1
X_07090_ _00892_ _00893_ _00894_ VPWR VGND _00895_ sg13g2_or3_1
X_07091_ _00883_ _00886_ _00891_ _00895_ VPWR VGND 
+ _00896_
+ sg13g2_nor4_2
X_07092_ _00896_ VPWR VGND _00897_ sg13g2_buf_8
X_07093_ \atbs_core_0.n1053_q\ VPWR VGND _00898_ sg13g2_inv_1
X_07094_ \atbs_core_0.spike_detector_0.lock_detection\ \atbs_core_0.detection_en\ \atbs_core_0.comp_upper_sync\ VPWR VGND _00899_ sg13g2_nand3b_1
X_07095_ _00898_ _00883_ _00899_ VPWR VGND _00900_ sg13g2_a21o_1
X_07096_ _00900_ VPWR VGND _00901_ sg13g2_buf_4
X_07097_ _00897_ _00901_ VPWR VGND _00902_ sg13g2_nor2_2
X_07098_ _00863_ _00882_ _00902_ VPWR VGND _00903_ sg13g2_a21oi_2
X_07099_ _00903_ VPWR VGND _00904_ sg13g2_buf_8
X_07100_ _00904_ VPWR VGND _00905_ sg13g2_buf_8
X_07101_ _00862_ _00905_ VPWR VGND _00906_ sg13g2_nand2_1
X_07102_ _00871_ VPWR VGND _00907_ sg13g2_inv_1
X_07103_ \atbs_core_0.adaptive_ctrl_0.delta_steps[0]\ VPWR VGND _00908_ sg13g2_buf_2
X_07104_ _00872_ VPWR VGND _00909_ sg13g2_inv_1
X_07105_ _00907_ \atbs_core_0.adaptive_ctrl_0.delta_steps[1]\ _00908_ _00909_ VPWR VGND 
+ _00910_
+ sg13g2_a22oi_1
X_07106_ \atbs_core_0.adaptive_ctrl_0.delta_steps[1]\ VPWR VGND _00911_ sg13g2_buf_2
X_07107_ \atbs_core_0.adaptive_ctrl_0.delta_steps[2]\ VPWR VGND _00912_ sg13g2_buf_2
X_07108_ _00912_ _00877_ VPWR VGND _00913_ sg13g2_nand2b_1
X_07109_ _00907_ _00911_ _00913_ VPWR VGND _00914_ sg13g2_o21ai_1
X_07110_ \atbs_core_0.adaptive_ctrl_0.delta_steps[3]\ VPWR VGND _00915_ sg13g2_buf_2
X_07111_ _00876_ _00915_ VPWR VGND _00916_ sg13g2_xor2_1
X_07112_ _00877_ \atbs_core_0.adaptive_ctrl_0.delta_steps[2]\ VPWR VGND _00917_ sg13g2_nor2b_1
X_07113_ \atbs_core_0.adaptive_ctrl_0.delta_steps[4]\ VPWR VGND _00918_ sg13g2_buf_4
X_07114_ _00869_ _00918_ VPWR VGND _00919_ sg13g2_nor2b_1
X_07115_ _00918_ _00869_ VPWR VGND _00920_ sg13g2_nor2b_1
X_07116_ _00916_ _00917_ _00919_ _00920_ VPWR VGND 
+ _00921_
+ sg13g2_nor4_1
X_07117_ _00910_ _00914_ _00921_ VPWR VGND _00922_ sg13g2_o21ai_1
X_07118_ _00876_ VPWR VGND _00923_ sg13g2_inv_1
X_07119_ _00923_ _00915_ _00919_ VPWR VGND _00924_ sg13g2_nor3_1
X_07120_ _00878_ VPWR VGND _00925_ sg13g2_inv_2
X_07121_ \atbs_core_0.adaptive_ctrl_0.delta_steps[7]\ VPWR VGND _00926_ sg13g2_buf_2
X_07122_ _00874_ VPWR VGND _00927_ sg13g2_inv_1
X_07123_ _00925_ _00926_ _00927_ VPWR VGND _00928_ sg13g2_o21ai_1
X_07124_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ _00868_ VPWR VGND _00929_ sg13g2_nand2b_1
X_07125_ \atbs_core_0.adaptive_ctrl_0.delta_steps[6]\ VPWR VGND _00930_ sg13g2_buf_4
X_07126_ _00930_ _00873_ VPWR VGND _00931_ sg13g2_nand2b_1
X_07127_ _00873_ _00930_ VPWR VGND _00932_ sg13g2_nor2b_1
X_07128_ _00929_ _00931_ _00932_ VPWR VGND _00933_ sg13g2_a21oi_1
X_07129_ _00920_ _00924_ _00928_ _00933_ VPWR VGND 
+ _00934_
+ sg13g2_nor4_2
X_07130_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ VPWR VGND _00935_ sg13g2_buf_4
X_07131_ _00868_ _00935_ VPWR VGND _00936_ sg13g2_nor2b_1
X_07132_ _00925_ _00926_ _00931_ _00936_ _00932_ VPWR 
+ VGND
+ _00937_ sg13g2_a221oi_1
X_07133_ _00928_ _00937_ VPWR VGND _00938_ sg13g2_nor2_1
X_07134_ _00922_ _00934_ _00938_ VPWR VGND _00939_ sg13g2_a21o_1
X_07135_ _00939_ VPWR VGND _00940_ sg13g2_buf_2
X_07136_ _00859_ _00023_ _00906_ _00940_ VPWR VGND 
+ _00941_
+ sg13g2_or4_1
X_07137_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ _00941_ VPWR VGND _00942_ sg13g2_and2_1
X_07138_ _00942_ VPWR VGND _00943_ sg13g2_buf_2
X_07139_ _00883_ VPWR VGND _00944_ sg13g2_buf_1
X_07140_ _00898_ _00944_ _00897_ VPWR VGND _00945_ sg13g2_a21oi_1
X_07141_ \atbs_core_0.comp_lower_sync\ _00867_ _00880_ VPWR VGND _00946_ sg13g2_nor3_1
X_07142_ \atbs_core_0.comp_upper_sync\ _00945_ _00946_ VPWR VGND _00947_ sg13g2_a21oi_1
X_07143_ _00864_ _00947_ VPWR VGND _00948_ sg13g2_or2_1
X_07144_ _00948_ VPWR VGND _00949_ sg13g2_buf_1
X_07145_ _00858_ _00949_ VPWR VGND _00950_ sg13g2_nor2_1
X_07146_ _00858_ _00943_ _00950_ VPWR VGND _00951_ sg13g2_a21oi_1
X_07147_ _00822_ _00824_ _00852_ _00951_ VPWR VGND 
+ _00952_
+ sg13g2_a22oi_1
X_07148_ _00952_ VPWR VGND \atbs_core_0.dac_control_0.dac_counter_strb\ sg13g2_buf_1
X_07149_ _00784_ VPWR VGND _00953_ sg13g2_inv_1
X_07150_ _00787_ _00953_ VPWR VGND _00954_ sg13g2_nand2_1
X_07151_ _00789_ _00785_ _00786_ VPWR VGND _00955_ sg13g2_nand3_1
X_07152_ \atbs_core_0.uart_0.uart_rx_0.n2873_o\ VPWR VGND _00956_ sg13g2_buf_1
X_07153_ _00753_ _00777_ VPWR VGND _00957_ sg13g2_or2_1
X_07154_ _00763_ _00753_ _00777_ VPWR VGND _00958_ sg13g2_nand3_1
X_07155_ _00763_ _00957_ _00958_ VPWR VGND _00959_ sg13g2_o21ai_1
X_07156_ _00759_ _00776_ VPWR VGND _00960_ sg13g2_xnor2_1
X_07157_ _00006_ _00959_ _00960_ VPWR VGND _00961_ sg13g2_nand3_1
X_07158_ _00773_ _00752_ VPWR VGND _00962_ sg13g2_or2_1
X_07159_ _00767_ _00773_ _00752_ VPWR VGND _00963_ sg13g2_nand3_1
X_07160_ _00767_ _00962_ _00963_ VPWR VGND _00964_ sg13g2_o21ai_1
X_07161_ _00771_ _00750_ VPWR VGND _00965_ sg13g2_xor2_1
X_07162_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ _00762_ VPWR VGND _00966_ sg13g2_xor2_1
X_07163_ _00755_ _00758_ VPWR VGND _00967_ sg13g2_xor2_1
X_07164_ _00965_ _00966_ _00967_ VPWR VGND _00968_ sg13g2_nor3_1
X_07165_ _00961_ _00964_ _00968_ VPWR VGND _00969_ sg13g2_nand3b_1
X_07166_ _00956_ _00969_ VPWR VGND _00970_ sg13g2_nand2_1
X_07167_ _00954_ _00955_ _00970_ VPWR VGND _00002_ sg13g2_o21ai_1
X_07168_ \atbs_core_0.uart_0.uart_rx_0.n2834_o\ VPWR VGND _00971_ sg13g2_buf_1
X_07169_ uart_rx_i VPWR VGND _00972_ sg13g2_inv_1
X_07170_ _00971_ _00972_ _00784_ _00748_ VPWR VGND 
+ _00973_
+ sg13g2_a22oi_1
X_07171_ _00973_ VPWR VGND _00001_ sg13g2_inv_1
X_07172_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[1]\ VPWR VGND _00974_ sg13g2_buf_1
X_07173_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[0]\ VPWR VGND _00975_ sg13g2_buf_1
X_07174_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[2]\ VPWR VGND _00976_ sg13g2_buf_1
X_07175_ _00974_ _00975_ _00976_ VPWR VGND _00977_ sg13g2_nand3_1
X_07176_ \atbs_core_0.uart_0.uart_tx_0.n2699_o\ VPWR VGND _00978_ sg13g2_buf_1
X_07177_ _00815_ _00977_ _00978_ VPWR VGND _00979_ sg13g2_o21ai_1
X_07178_ _00792_ _00815_ _00979_ VPWR VGND _00005_ sg13g2_o21ai_1
X_07179_ _00818_ _00031_ VPWR VGND _00980_ sg13g2_nor2_1
X_07180_ _00816_ _00980_ _00815_ VPWR VGND _00981_ sg13g2_o21ai_1
X_07181_ _00981_ VPWR VGND _00004_ sg13g2_inv_1
X_07182_ \atbs_core_0.enable_read\ VPWR VGND _00982_ sg13g2_inv_1
X_07183_ \atbs_core_0.spike_memory_0.head[1]\ \atbs_core_0.spike_memory_0.n1973_q[1]\ VPWR VGND _00983_ sg13g2_xor2_1
X_07184_ _00983_ VPWR VGND _00984_ sg13g2_buf_1
X_07185_ \atbs_core_0.spike_memory_0.n1973_q[0]\ VPWR VGND _00985_ sg13g2_buf_1
X_07186_ \atbs_core_0.spike_memory_0.head[0]\ VPWR VGND _00986_ sg13g2_buf_1
X_07187_ _00985_ _00986_ VPWR VGND _00987_ sg13g2_nor2b_1
X_07188_ _00986_ _00985_ VPWR VGND _00988_ sg13g2_nor2b_1
X_07189_ _00984_ _00987_ _00988_ VPWR VGND _00989_ sg13g2_nor3_1
X_07190_ _00982_ \atbs_core_0.spike_memory_0.n1912_o\ _00989_ VPWR VGND _00990_ sg13g2_nor3_1
X_07191_ _00990_ VPWR VGND \atbs_core_0.spike_memory_0.n1914_o\ sg13g2_buf_1
X_07192_ \atbs_core_0.spike_detector_0.n1258_q\ \atbs_core_0.spike_detector_0.lower_is_changing\ VPWR VGND _00991_ sg13g2_nor2_1
X_07193_ _00991_ VPWR VGND \atbs_core_0.spike_detector_0.n1246_o\ sg13g2_inv_1
X_07194_ _00904_ VPWR VGND _00992_ sg13g2_inv_16
X_07195_ _00935_ VPWR VGND _00993_ sg13g2_inv_1
X_07196_ _00930_ _00890_ VPWR VGND _00994_ sg13g2_nor2b_1
X_07197_ _00889_ _00918_ VPWR VGND _00995_ sg13g2_nand2b_1
X_07198_ _00993_ _00994_ _00995_ VPWR VGND _00996_ sg13g2_nor3_1
X_07199_ _00930_ VPWR VGND _00997_ sg13g2_inv_1
X_07200_ _00890_ _00997_ _00993_ _00995_ _00888_ VPWR 
+ VGND
+ _00998_ sg13g2_a221oi_1
X_07201_ _00890_ _00997_ _00026_ VPWR VGND _00999_ sg13g2_o21ai_1
X_07202_ _00996_ _00998_ _00999_ VPWR VGND _01000_ sg13g2_or3_1
X_07203_ _00884_ _00885_ VPWR VGND _01001_ sg13g2_nor2_1
X_07204_ _00926_ _01000_ _01001_ VPWR VGND _01002_ sg13g2_o21ai_1
X_07205_ _01002_ VPWR VGND _01003_ sg13g2_buf_2
X_07206_ _00892_ _00908_ VPWR VGND _01004_ sg13g2_nor2b_1
X_07207_ _00911_ _01004_ VPWR VGND _01005_ sg13g2_nor2_1
X_07208_ _00893_ VPWR VGND _01006_ sg13g2_inv_1
X_07209_ _00894_ _00912_ VPWR VGND _01007_ sg13g2_nor2b_1
X_07210_ _01006_ _00915_ _00911_ _01004_ _01007_ VPWR 
+ VGND
+ _01008_ sg13g2_a221oi_1
X_07211_ _00887_ _01005_ _01008_ VPWR VGND _01009_ sg13g2_o21ai_1
X_07212_ _00915_ VPWR VGND _01010_ sg13g2_inv_1
X_07213_ _00912_ _00894_ VPWR VGND _01011_ sg13g2_nor2b_1
X_07214_ _01010_ _01011_ _00893_ VPWR VGND _01012_ sg13g2_o21ai_1
X_07215_ _00918_ VPWR VGND _01013_ sg13g2_inv_1
X_07216_ _00915_ _00912_ VPWR VGND _01014_ sg13g2_nor2_1
X_07217_ _00889_ _01013_ _01014_ _00894_ _00885_ VPWR 
+ VGND
+ _01015_ sg13g2_a221oi_1
X_07218_ _00926_ VPWR VGND _01016_ sg13g2_inv_1
X_07219_ _00884_ _01016_ _00993_ _00888_ _00994_ VPWR 
+ VGND
+ _01017_ sg13g2_a221oi_1
X_07220_ _01012_ _01015_ _01017_ VPWR VGND _01018_ sg13g2_and3_1
X_07221_ _00885_ _00926_ VPWR VGND _01019_ sg13g2_nor2b_1
X_07222_ _01009_ _01018_ _01000_ _01019_ VPWR VGND 
+ _01020_
+ sg13g2_a22oi_1
X_07223_ _01020_ VPWR VGND _01021_ sg13g2_buf_4
X_07224_ _00992_ _01003_ _01021_ VPWR VGND _01022_ sg13g2_and3_2
X_07225_ _01022_ VPWR VGND _01023_ sg13g2_buf_8
X_07226_ _00860_ _01023_ VPWR VGND _01024_ sg13g2_nor2_1
X_07227_ _00992_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.spike_i\ sg13g2_buf_8
X_07228_ _00029_ \atbs_core_0.adaptive_ctrl_0.spike_i\ VPWR VGND _01025_ sg13g2_nand2_1
X_07229_ _01025_ VPWR VGND _01026_ sg13g2_buf_2
X_07230_ _00859_ _00023_ _01024_ _01026_ VPWR VGND 
+ _01027_
+ sg13g2_nor4_1
X_07231_ _01027_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ VPWR VGND _01028_ sg13g2_nand2b_1
X_07232_ _01028_ VPWR VGND _01029_ sg13g2_buf_1
X_07233_ _01029_ VPWR VGND _01030_ sg13g2_inv_1
X_07234_ _00858_ _01030_ _00950_ VPWR VGND _01031_ sg13g2_a21oi_1
X_07235_ _00852_ _01031_ VPWR VGND _01032_ sg13g2_nand2_1
X_07236_ _00853_ \atbs_core_0.debouncer_4.debounced\ VPWR VGND _01033_ sg13g2_nor2b_1
X_07237_ _00853_ \atbs_core_0.enable_analog_uart\ _01033_ VPWR VGND _01034_ sg13g2_a21o_1
X_07238_ _01034_ VPWR VGND _01035_ sg13g2_buf_1
X_07239_ _01032_ _01035_ \atbs_core_0.dac_control_1.n1629_o\ VPWR VGND \atbs_core_0.dac_control_1.n1632_o\ sg13g2_mux2_1
X_07240_ \atbs_core_0.dac_control_1.n1721_q\ VPWR VGND _01036_ sg13g2_buf_4
X_07241_ _01036_ VPWR VGND _01037_ sg13g2_inv_1
X_07242_ _00852_ _01031_ VPWR VGND _01038_ sg13g2_and2_1
X_07243_ _01038_ VPWR VGND _01039_ sg13g2_buf_1
X_07244_ \atbs_core_0.dac_control_1.n1629_o\ _01037_ _01039_ VPWR VGND \atbs_core_0.dac_control_1.dac_counter_strb\ sg13g2_a21oi_1
X_07245_ _00978_ VPWR VGND _01040_ sg13g2_inv_1
X_07246_ _01040_ _00977_ VPWR VGND _01041_ sg13g2_nor2_1
X_07247_ _01041_ \atbs_core_0.uart_0.uart_tx_0.n2758_o\ _00815_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2766_o[2]\ sg13g2_mux2_1
X_07248_ \atbs_core_0.uart_0.rx_data_strb_o\ VPWR VGND _01042_ sg13g2_inv_1
X_07249_ _01042_ \atbs_core_0.n1061_q\ \atbs_core_0.analog_trigger_uart\ VPWR VGND _01043_ sg13g2_nor3_1
X_07250_ \atbs_core_0.uart_0.uart_rx_0.n2915_o\ VPWR VGND _01044_ sg13g2_inv_1
X_07251_ \atbs_core_0.uart_0.uart_rx_0.n2921_o\ \atbs_core_0.uart_0.uart_rx_0.n2919_o\ VPWR VGND _01045_ sg13g2_nand2b_1
X_07252_ \atbs_core_0.uart_0.uart_rx_0.n2917_o\ _01044_ _01045_ VPWR VGND _01046_ sg13g2_nor3_1
X_07253_ _00049_ _01046_ VPWR VGND _01047_ sg13g2_nand2_1
X_07254_ \atbs_core_0.uart_0.uart_rx_0.n2907_o\ VPWR VGND _01048_ sg13g2_buf_1
X_07255_ \atbs_core_0.atbs_win_length_uart\ VPWR VGND _01049_ sg13g2_buf_1
X_07256_ _01049_ \atbs_core_0.atbs_max_delta_steps_uart\ VPWR VGND _01050_ sg13g2_nor2_1
X_07257_ \atbs_core_0.uart_0.uart_rx_0.n2909_o\ VPWR VGND _01051_ sg13g2_buf_1
X_07258_ \atbs_core_0.uart_0.uart_rx_0.n2913_o\ VPWR VGND _01052_ sg13g2_buf_1
X_07259_ \atbs_core_0.uart_0.uart_rx_0.n2911_o\ VPWR VGND _01053_ sg13g2_buf_1
X_07260_ _01052_ _01053_ VPWR VGND _01054_ sg13g2_nor2b_1
X_07261_ _01051_ _01054_ VPWR VGND _01055_ sg13g2_nor2b_1
X_07262_ \atbs_core_0.uart_0.uart_rx_0.n2917_o\ VPWR VGND _01056_ sg13g2_inv_1
X_07263_ _01056_ _01044_ \atbs_core_0.uart_0.uart_rx_0.n2921_o\ \atbs_core_0.uart_0.uart_rx_0.n2919_o\ VPWR VGND 
+ _01057_
+ sg13g2_or4_1
X_07264_ _01057_ VPWR VGND _01058_ sg13g2_buf_1
X_07265_ _01048_ _01050_ _01055_ _01058_ VPWR VGND 
+ _01059_
+ sg13g2_nand4_1
X_07266_ _01047_ _01059_ _00048_ VPWR VGND _01060_ sg13g2_o21ai_1
X_07267_ \atbs_core_0.debouncer_5.debounced\ \atbs_core_0.n1049_q\ VPWR VGND _01061_ sg13g2_xor2_1
X_07268_ \atbs_core_0.adaptive_mode_d\ \atbs_core_0.adaptive_mode_debounced\ VPWR VGND _01062_ sg13g2_xor2_1
X_07269_ _00853_ \atbs_core_0.control_mode_d\ VPWR VGND _01063_ sg13g2_xor2_1
X_07270_ _01061_ _01062_ _01063_ VPWR VGND _01064_ sg13g2_nor3_1
X_07271_ \atbs_core_0.n1050_q\ \atbs_core_0.debouncer_0.debounced\ VPWR VGND _01065_ sg13g2_xnor2_1
X_07272_ \atbs_core_0.n1048_q\ \atbs_core_0.debouncer_3.debounced\ VPWR VGND _01066_ sg13g2_xnor2_1
X_07273_ _01064_ _01065_ _01066_ VPWR VGND _01067_ sg13g2_nand3_1
X_07274_ _01043_ _01060_ _01067_ VPWR VGND _01068_ sg13g2_a21oi_1
X_07275_ _00849_ VPWR VGND _01069_ sg13g2_buf_1
X_07276_ _01069_ _00843_ VPWR VGND _01070_ sg13g2_nor2_1
X_07277_ _00849_ VPWR VGND _01071_ sg13g2_inv_1
X_07278_ _01071_ _00844_ VPWR VGND _01072_ sg13g2_nor2_1
X_07279_ _01070_ _01072_ _00842_ VPWR VGND _01073_ sg13g2_o21ai_1
X_07280_ _01068_ _01073_ VPWR VGND _01074_ sg13g2_nor2_1
X_07281_ \atbs_core_0.atbs_max_delta_steps_uart\ VPWR VGND _01075_ sg13g2_inv_1
X_07282_ \atbs_core_0.n1067_q\ VPWR VGND _01076_ sg13g2_inv_1
X_07283_ \atbs_core_0.baudrate_uart\ VPWR VGND _01077_ sg13g2_buf_1
X_07284_ _01077_ _01043_ VPWR VGND _01078_ sg13g2_nor2b_1
X_07285_ _01076_ _01078_ VPWR VGND _01079_ sg13g2_and2_1
X_07286_ _01079_ VPWR VGND _01080_ sg13g2_buf_1
X_07287_ _01049_ _01080_ VPWR VGND _01081_ sg13g2_nor2b_1
X_07288_ _01053_ _01052_ VPWR VGND _01082_ sg13g2_nor2_1
X_07289_ _01051_ _01082_ VPWR VGND _01083_ sg13g2_nand2_1
X_07290_ _01048_ _01083_ VPWR VGND _01084_ sg13g2_nor2_1
X_07291_ _01075_ _01081_ _01046_ _01084_ VPWR VGND 
+ _01085_
+ sg13g2_nand4_1
X_07292_ \atbs_core_0.n31_o\ _01085_ VPWR VGND _00120_ sg13g2_and2_1
X_07293_ _01074_ _00120_ VPWR VGND _00119_ sg13g2_nor2b_1
X_07294_ \atbs_core_0.debouncer_0.debounced\ \atbs_core_0.n1078_q\ _00853_ VPWR VGND _01086_ sg13g2_mux2_1
X_07295_ _01048_ VPWR VGND _01087_ sg13g2_inv_1
X_07296_ _01087_ _01083_ VPWR VGND _01088_ sg13g2_nor2_1
X_07297_ _01080_ _01046_ _01050_ _01088_ VPWR VGND 
+ _01089_
+ sg13g2_nand4_1
X_07298_ \atbs_core_0.n1051_q\ \atbs_core_0.n37_o\ VPWR VGND _01090_ sg13g2_nand2b_1
X_07299_ _01086_ _01089_ _01090_ VPWR VGND _01091_ sg13g2_and3_1
X_07300_ _01091_ VPWR VGND _01092_ sg13g2_buf_1
X_07301_ _00849_ _00842_ VPWR VGND _01093_ sg13g2_nand2_1
X_07302_ _00843_ _01092_ _01093_ VPWR VGND _01094_ sg13g2_nor3_1
X_07303_ _01094_ VPWR VGND _01095_ sg13g2_buf_1
X_07304_ _01086_ _01095_ VPWR VGND _01096_ sg13g2_nand2_1
X_07305_ _00119_ _01096_ VPWR VGND _00122_ sg13g2_and2_1
X_07306_ \atbs_core_0.adaptive_ctrl_0.n1308_o\ VPWR VGND _01097_ sg13g2_buf_1
X_07307_ _00911_ VPWR VGND _01098_ sg13g2_inv_1
X_07308_ _01013_ _01098_ _01014_ VPWR VGND _01099_ sg13g2_nand3_1
X_07309_ _00926_ _00930_ _00935_ _01099_ VPWR VGND 
+ _01100_
+ sg13g2_nor4_1
X_07310_ _00908_ _01100_ VPWR VGND _01101_ sg13g2_nand2_1
X_07311_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _01097_ _01101_ VPWR VGND _01102_ sg13g2_nand3_1
X_07312_ _00862_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ _01102_ VPWR VGND _00125_ sg13g2_o21ai_1
X_07313_ _00052_ VPWR VGND _01103_ sg13g2_buf_1
X_07314_ _01103_ VPWR VGND _01104_ sg13g2_inv_1
X_07315_ _00949_ VPWR VGND _01105_ sg13g2_inv_1
X_07316_ _01105_ VPWR VGND _01106_ sg13g2_buf_1
X_07317_ _01106_ VPWR VGND _01107_ sg13g2_buf_1
X_07318_ _01104_ _01107_ VPWR VGND _01108_ sg13g2_nor2_1
X_07319_ _01097_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _01108_ VPWR VGND _00126_ sg13g2_mux2_1
X_07320_ \atbs_core_0.adaptive_ctrl_0.n1447_q[0]\ VPWR VGND _01109_ sg13g2_buf_1
X_07321_ _01109_ VPWR VGND _01110_ sg13g2_inv_1
X_07322_ \atbs_core_0.adaptive_ctrl_0.adaptive_strb\ _00905_ _00940_ VPWR VGND _01111_ sg13g2_nand3_1
X_07323_ _01003_ _01021_ _00904_ VPWR VGND _01112_ sg13g2_a21o_1
X_07324_ _00859_ _01112_ VPWR VGND _01113_ sg13g2_or2_1
X_07325_ _00029_ VPWR VGND _01114_ sg13g2_inv_1
X_07326_ _01111_ _01113_ _01114_ VPWR VGND _01115_ sg13g2_a21oi_1
X_07327_ _01115_ VPWR VGND _01116_ sg13g2_buf_1
X_07328_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[2]\ VPWR VGND _01117_ sg13g2_a21oi_1
X_07329_ _00997_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[6]\ _00032_ VPWR VGND _01118_ sg13g2_o21ai_1
X_07330_ _01013_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ VPWR VGND _01119_ sg13g2_nand2_1
X_07331_ _00912_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ VPWR VGND _01120_ sg13g2_nor2b_1
X_07332_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _01120_ VPWR VGND _01121_ sg13g2_nand2_1
X_07333_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _01120_ _01010_ VPWR VGND _01122_ sg13g2_o21ai_1
X_07334_ _01119_ _01121_ _01122_ VPWR VGND _01123_ sg13g2_nand3_1
X_07335_ _01013_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _01123_ VPWR VGND _01124_ sg13g2_o21ai_1
X_07336_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[5]\ VPWR VGND _01125_ sg13g2_inv_1
X_07337_ _00935_ _01124_ _01125_ VPWR VGND _01126_ sg13g2_o21ai_1
X_07338_ _00935_ _01124_ VPWR VGND _01127_ sg13g2_nand2_1
X_07339_ _00997_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[6]\ _01126_ _01127_ VPWR VGND 
+ _01128_
+ sg13g2_a22oi_1
X_07340_ _01117_ _01118_ _01128_ VPWR VGND _01129_ sg13g2_nor3_1
X_07341_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[2]\ _01100_ VPWR VGND _01130_ sg13g2_nor3_1
X_07342_ \atbs_core_0.adaptive_ctrl_0.n1352_o\ VPWR VGND _01131_ sg13g2_buf_1
X_07343_ _01129_ _01130_ _01131_ VPWR VGND _01132_ sg13g2_o21ai_1
X_07344_ _01132_ VPWR VGND _01133_ sg13g2_buf_1
X_07345_ _01129_ VPWR VGND _01134_ sg13g2_inv_1
X_07346_ _00911_ _01134_ _01133_ VPWR VGND _01135_ sg13g2_a21oi_1
X_07347_ _00090_ _01133_ _01135_ VPWR VGND _01136_ sg13g2_a21oi_1
X_07348_ _01095_ _01116_ _01136_ VPWR VGND _01137_ sg13g2_nor3_1
X_07349_ _01110_ _01116_ _01137_ VPWR VGND _00127_ sg13g2_a21o_1
X_07350_ _01133_ VPWR VGND _01138_ sg13g2_buf_1
X_07351_ _01129_ VPWR VGND _01139_ sg13g2_buf_1
X_07352_ _00043_ _01139_ VPWR VGND _01140_ sg13g2_nor2_1
X_07353_ _00908_ _01139_ _01140_ VPWR VGND _01141_ sg13g2_a21oi_1
X_07354_ _01133_ _01141_ VPWR VGND _01142_ sg13g2_nor2_1
X_07355_ _00911_ _01138_ _01142_ VPWR VGND _01143_ sg13g2_a21oi_1
X_07356_ _01095_ _01115_ VPWR VGND _01144_ sg13g2_or2_1
X_07357_ _01144_ VPWR VGND _01145_ sg13g2_buf_1
X_07358_ \atbs_core_0.adaptive_ctrl_0.n1447_q[1]\ VPWR VGND _01146_ sg13g2_buf_1
X_07359_ _01146_ _01116_ VPWR VGND _01147_ sg13g2_nand2_1
X_07360_ _01143_ _01145_ _01147_ VPWR VGND _00128_ sg13g2_o21ai_1
X_07361_ _00045_ VPWR VGND _01148_ sg13g2_inv_1
X_07362_ _00040_ _01139_ VPWR VGND _01149_ sg13g2_nor2_1
X_07363_ _01148_ _01139_ _01149_ VPWR VGND _01150_ sg13g2_a21oi_1
X_07364_ _01138_ _01150_ VPWR VGND _01151_ sg13g2_nor2_1
X_07365_ _00912_ _01138_ _01151_ VPWR VGND _01152_ sg13g2_a21oi_1
X_07366_ \atbs_core_0.adaptive_ctrl_0.n1447_q[2]\ VPWR VGND _01153_ sg13g2_buf_1
X_07367_ _01153_ _01116_ VPWR VGND _01154_ sg13g2_nand2_1
X_07368_ _01145_ _01152_ _01154_ VPWR VGND _00129_ sg13g2_o21ai_1
X_07369_ _00043_ VPWR VGND _01155_ sg13g2_inv_1
X_07370_ _00039_ _01139_ VPWR VGND _01156_ sg13g2_nor2_1
X_07371_ _01155_ _01139_ _01156_ VPWR VGND _01157_ sg13g2_a21oi_1
X_07372_ _01138_ _01157_ VPWR VGND _01158_ sg13g2_nor2_1
X_07373_ _00915_ _01138_ _01158_ VPWR VGND _01159_ sg13g2_a21oi_1
X_07374_ \atbs_core_0.adaptive_ctrl_0.n1447_q[3]\ _01116_ VPWR VGND _01160_ sg13g2_nand2_1
X_07375_ _01145_ _01159_ _01160_ VPWR VGND _00130_ sg13g2_o21ai_1
X_07376_ _00040_ VPWR VGND _01161_ sg13g2_inv_1
X_07377_ _00036_ _01139_ VPWR VGND _01162_ sg13g2_nor2_1
X_07378_ _01161_ _01139_ _01162_ VPWR VGND _01163_ sg13g2_a21oi_1
X_07379_ _01138_ _01163_ VPWR VGND _01164_ sg13g2_nor2_1
X_07380_ _00918_ _01138_ _01164_ VPWR VGND _01165_ sg13g2_a21oi_1
X_07381_ \atbs_core_0.adaptive_ctrl_0.n1447_q[4]\ VPWR VGND _01166_ sg13g2_buf_1
X_07382_ _01166_ _01116_ VPWR VGND _01167_ sg13g2_nand2_1
X_07383_ _01145_ _01165_ _01167_ VPWR VGND _00131_ sg13g2_o21ai_1
X_07384_ _00035_ VPWR VGND _01168_ sg13g2_inv_1
X_07385_ _00039_ _01139_ VPWR VGND _01169_ sg13g2_nand2_1
X_07386_ _01168_ _01139_ _01169_ VPWR VGND _01170_ sg13g2_o21ai_1
X_07387_ _01133_ _01170_ VPWR VGND _01171_ sg13g2_nor2_1
X_07388_ _00935_ _01138_ _01171_ VPWR VGND _01172_ sg13g2_a21oi_1
X_07389_ \atbs_core_0.adaptive_ctrl_0.n1447_q[5]\ VPWR VGND _01173_ sg13g2_buf_1
X_07390_ _01173_ _01116_ VPWR VGND _01174_ sg13g2_nand2_1
X_07391_ _01145_ _01172_ _01174_ VPWR VGND _00132_ sg13g2_o21ai_1
X_07392_ \atbs_core_0.adaptive_ctrl_0.n1447_q[6]\ VPWR VGND _01175_ sg13g2_buf_1
X_07393_ _00036_ _01129_ VPWR VGND _01176_ sg13g2_nand2b_1
X_07394_ _00032_ _01176_ _01133_ VPWR VGND _01177_ sg13g2_a21oi_1
X_07395_ _00930_ _01133_ _01177_ VPWR VGND _01178_ sg13g2_a21oi_1
X_07396_ _01095_ _01116_ _01178_ VPWR VGND _01179_ sg13g2_nor3_1
X_07397_ _01175_ _01116_ _01179_ VPWR VGND _00133_ sg13g2_a21o_1
X_07398_ _00997_ _01134_ _01133_ VPWR VGND _01180_ sg13g2_nor3_1
X_07399_ _00926_ _01138_ _01180_ VPWR VGND _01181_ sg13g2_a21oi_1
X_07400_ \atbs_core_0.adaptive_ctrl_0.n1447_q[7]\ _01116_ VPWR VGND _01182_ sg13g2_nand2_1
X_07401_ _01145_ _01181_ _01182_ VPWR VGND _00134_ sg13g2_o21ai_1
X_07402_ _00843_ _01092_ VPWR VGND _01183_ sg13g2_nor2_1
X_07403_ _01093_ _01183_ VPWR VGND _01184_ sg13g2_nand2b_1
X_07404_ _01184_ VPWR VGND _01185_ sg13g2_buf_1
X_07405_ _01131_ VPWR VGND _01186_ sg13g2_buf_1
X_07406_ _00908_ _01131_ VPWR VGND _01187_ sg13g2_nand2_1
X_07407_ _01186_ _00091_ _01187_ VPWR VGND _01188_ sg13g2_o21ai_1
X_07408_ _01185_ _01188_ VPWR VGND _00135_ sg13g2_nand2_1
X_07409_ _01095_ VPWR VGND _01189_ sg13g2_buf_1
X_07410_ _01186_ _01146_ VPWR VGND _01190_ sg13g2_nor2b_1
X_07411_ _00911_ _01186_ _01190_ VPWR VGND _01191_ sg13g2_a21oi_1
X_07412_ _01189_ _01191_ VPWR VGND _00136_ sg13g2_nor2_1
X_07413_ _01186_ _01153_ VPWR VGND _01192_ sg13g2_nor2b_1
X_07414_ _00912_ _01186_ _01192_ VPWR VGND _01193_ sg13g2_a21oi_1
X_07415_ _01189_ _01193_ VPWR VGND _00137_ sg13g2_nor2_1
X_07416_ \atbs_core_0.adaptive_ctrl_0.n1447_q[3]\ VPWR VGND _01194_ sg13g2_inv_1
X_07417_ _01194_ _01010_ _01186_ VPWR VGND _01195_ sg13g2_mux2_1
X_07418_ _01189_ _01195_ VPWR VGND _00138_ sg13g2_nor2_1
X_07419_ _01131_ _01166_ VPWR VGND _01196_ sg13g2_nor2b_1
X_07420_ _00918_ _01186_ _01196_ VPWR VGND _01197_ sg13g2_a21oi_1
X_07421_ _01189_ _01197_ VPWR VGND _00139_ sg13g2_nor2_1
X_07422_ _01131_ _01173_ VPWR VGND _01198_ sg13g2_nor2b_1
X_07423_ _00935_ _01186_ _01198_ VPWR VGND _01199_ sg13g2_a21oi_1
X_07424_ _01189_ _01199_ VPWR VGND _00140_ sg13g2_nor2_1
X_07425_ _01131_ _01175_ VPWR VGND _01200_ sg13g2_nor2b_1
X_07426_ _00930_ _01186_ _01200_ VPWR VGND _01201_ sg13g2_a21oi_1
X_07427_ _01189_ _01201_ VPWR VGND _00141_ sg13g2_nor2_1
X_07428_ _01131_ \atbs_core_0.adaptive_ctrl_0.n1447_q[7]\ VPWR VGND _01202_ sg13g2_nor2b_1
X_07429_ _00926_ _01186_ _01202_ VPWR VGND _01203_ sg13g2_a21oi_1
X_07430_ _01189_ _01203_ VPWR VGND _00142_ sg13g2_nor2_1
X_07431_ _00943_ VPWR VGND _01204_ sg13g2_buf_1
X_07432_ _01204_ _00092_ VPWR VGND _01205_ sg13g2_nand2b_1
X_07433_ _00859_ _00860_ \atbs_core_0.adaptive_ctrl_0.n1444_q\ VPWR VGND _01206_ sg13g2_nor3_1
X_07434_ _00928_ _00937_ _01206_ VPWR VGND _01207_ sg13g2_o21ai_1
X_07435_ _00922_ _00934_ _01207_ VPWR VGND _01208_ sg13g2_a21oi_1
X_07436_ _01208_ VPWR VGND _01209_ sg13g2_buf_2
X_07437_ _00905_ _01209_ VPWR VGND _01210_ sg13g2_nand2_2
X_07438_ _01210_ VPWR VGND _01211_ sg13g2_buf_4
X_07439_ _00908_ VPWR VGND _01212_ sg13g2_inv_1
X_07440_ _00904_ _00940_ _01212_ VPWR VGND _01213_ sg13g2_a21oi_1
X_07441_ _00892_ _00992_ VPWR VGND _01214_ sg13g2_and2_1
X_07442_ _01003_ VPWR VGND _01215_ sg13g2_buf_4
X_07443_ _01021_ VPWR VGND _01216_ sg13g2_buf_4
X_07444_ _01215_ _01216_ VPWR VGND _01217_ sg13g2_nand2_1
X_07445_ _00922_ _00934_ _00938_ VPWR VGND _01218_ sg13g2_a21oi_1
X_07446_ _01218_ VPWR VGND _01219_ sg13g2_buf_4
X_07447_ _00897_ _00901_ _00872_ VPWR VGND _01220_ sg13g2_o21ai_1
X_07448_ _00863_ _00882_ _01220_ VPWR VGND _01221_ sg13g2_a21o_1
X_07449_ _01219_ _01221_ _00861_ VPWR VGND _01222_ sg13g2_o21ai_1
X_07450_ _01112_ _01213_ _01214_ _01217_ _01222_ VPWR 
+ VGND
+ _01223_ sg13g2_a221oi_1
X_07451_ _01223_ VPWR VGND _01224_ sg13g2_buf_2
X_07452_ _01212_ _01110_ _01206_ VPWR VGND _01225_ sg13g2_and3_1
X_07453_ _00897_ _00901_ _01225_ VPWR VGND _01226_ sg13g2_o21ai_1
X_07454_ _00863_ _00882_ _01226_ VPWR VGND _01227_ sg13g2_a21oi_1
X_07455_ _00908_ _00862_ VPWR VGND _01228_ sg13g2_nor2_1
X_07456_ _01219_ _01227_ _01228_ VPWR VGND _01229_ sg13g2_a21oi_1
X_07457_ _00908_ _01109_ VPWR VGND _01230_ sg13g2_nand2_1
X_07458_ _01230_ VPWR VGND _01231_ sg13g2_inv_1
X_07459_ _00905_ _01209_ _01231_ VPWR VGND _01232_ sg13g2_nand3_1
X_07460_ _01229_ _01232_ VPWR VGND _01233_ sg13g2_nand2_1
X_07461_ _01211_ _01224_ _01233_ VPWR VGND _01234_ sg13g2_a21oi_1
X_07462_ _01234_ VPWR VGND _01235_ sg13g2_buf_2
X_07463_ _00892_ _01235_ VPWR VGND _01236_ sg13g2_xnor2_1
X_07464_ _01204_ _01236_ VPWR VGND _01237_ sg13g2_nand2_1
X_07465_ _01095_ VPWR VGND _01238_ sg13g2_buf_1
X_07466_ _01205_ _01237_ _01238_ VPWR VGND _00143_ sg13g2_a21oi_1
X_07467_ _00892_ _01026_ VPWR VGND _01239_ sg13g2_xnor2_1
X_07468_ _01235_ _01239_ VPWR VGND _01240_ sg13g2_nand2_1
X_07469_ _00046_ VPWR VGND _01241_ sg13g2_inv_1
X_07470_ _00897_ _00901_ VPWR VGND _01242_ sg13g2_or2_1
X_07471_ _01242_ VPWR VGND _01243_ sg13g2_buf_2
X_07472_ _01243_ VPWR VGND _01244_ sg13g2_buf_4
X_07473_ _00863_ _00882_ VPWR VGND _01245_ sg13g2_nand2_1
X_07474_ _01245_ VPWR VGND _01246_ sg13g2_buf_4
X_07475_ _00860_ _00045_ VPWR VGND _01247_ sg13g2_nand2_1
X_07476_ _01241_ _01247_ VPWR VGND _01248_ sg13g2_nand2_1
X_07477_ _01244_ _01246_ _01215_ _01216_ _01248_ VPWR 
+ VGND
+ _01249_ sg13g2_a221oi_1
X_07478_ _00904_ _01209_ _01148_ VPWR VGND _01250_ sg13g2_a21oi_1
X_07479_ _00871_ _00904_ _00940_ _01247_ VPWR VGND 
+ _01251_
+ sg13g2_nand4_1
X_07480_ _01249_ _01250_ _01251_ VPWR VGND _01252_ sg13g2_nand3b_1
X_07481_ _01252_ VPWR VGND _01253_ sg13g2_buf_4
X_07482_ _00871_ _00992_ _01219_ VPWR VGND _01254_ sg13g2_nor3_1
X_07483_ _01243_ _01246_ _01003_ _01021_ _01241_ VPWR 
+ VGND
+ _01255_ sg13g2_a221oi_1
X_07484_ _00905_ _01209_ _00860_ VPWR VGND _01256_ sg13g2_a21oi_1
X_07485_ _01254_ _01255_ _01256_ VPWR VGND _01257_ sg13g2_o21ai_1
X_07486_ _01257_ VPWR VGND _01258_ sg13g2_buf_2
X_07487_ _00904_ _01209_ VPWR VGND _01259_ sg13g2_and2_1
X_07488_ _01259_ VPWR VGND _01260_ sg13g2_buf_2
X_07489_ _00911_ _01146_ VPWR VGND _01261_ sg13g2_xnor2_1
X_07490_ _01230_ _01261_ VPWR VGND _01262_ sg13g2_xnor2_1
X_07491_ _01260_ _01262_ VPWR VGND _01263_ sg13g2_nand2_1
X_07492_ _01253_ _01258_ _01263_ VPWR VGND _01264_ sg13g2_and3_1
X_07493_ _01264_ VPWR VGND _01265_ sg13g2_buf_1
X_07494_ _01241_ _01265_ VPWR VGND _01266_ sg13g2_xnor2_1
X_07495_ _01240_ _01266_ VPWR VGND _01267_ sg13g2_xnor2_1
X_07496_ _00943_ _01267_ VPWR VGND _01268_ sg13g2_nand2_1
X_07497_ _00887_ _01204_ _01268_ VPWR VGND _01269_ sg13g2_o21ai_1
X_07498_ _01189_ _01269_ VPWR VGND _00144_ sg13g2_nor2_1
X_07499_ _01241_ _01026_ _01265_ VPWR VGND _01270_ sg13g2_nand3_1
X_07500_ _00887_ _01235_ VPWR VGND _01271_ sg13g2_nand2b_1
X_07501_ _00892_ _01270_ _01271_ VPWR VGND _01272_ sg13g2_a21oi_1
X_07502_ _01253_ _01258_ _01026_ VPWR VGND _01273_ sg13g2_a21o_1
X_07503_ _01114_ _00905_ VPWR VGND _01274_ sg13g2_nor2_1
X_07504_ _01241_ _01274_ _00892_ VPWR VGND _01275_ sg13g2_o21ai_1
X_07505_ _01235_ _01273_ _01275_ VPWR VGND _01276_ sg13g2_nand3_1
X_07506_ _00887_ _00046_ VPWR VGND _01277_ sg13g2_or2_1
X_07507_ _01277_ _01241_ _01265_ VPWR VGND _01278_ sg13g2_mux2_1
X_07508_ _00892_ _01241_ _01265_ VPWR VGND _01279_ sg13g2_a21o_1
X_07509_ _01026_ _01235_ VPWR VGND _01280_ sg13g2_and2_1
X_07510_ _01276_ _01278_ _01279_ _01280_ VPWR VGND 
+ _01281_
+ sg13g2_a22oi_1
X_07511_ _01272_ _01281_ VPWR VGND _01282_ sg13g2_nor2_1
X_07512_ _00912_ _01153_ VPWR VGND _01283_ sg13g2_xor2_1
X_07513_ _00908_ _01109_ _01146_ VPWR VGND _01284_ sg13g2_a21o_1
X_07514_ _00908_ _01146_ _01109_ VPWR VGND _01285_ sg13g2_and3_1
X_07515_ _00911_ _01284_ _01285_ VPWR VGND _01286_ sg13g2_a21oi_1
X_07516_ _01283_ _01286_ VPWR VGND _01287_ sg13g2_xnor2_1
X_07517_ _01210_ _01287_ VPWR VGND _01288_ sg13g2_nor2_1
X_07518_ _00877_ VPWR VGND _01289_ sg13g2_inv_1
X_07519_ _01289_ _00860_ VPWR VGND _01290_ sg13g2_nor2_1
X_07520_ _00897_ _00901_ _01290_ VPWR VGND _01291_ sg13g2_o21ai_1
X_07521_ _00863_ _00882_ _01291_ VPWR VGND _01292_ sg13g2_a21oi_1
X_07522_ _00897_ _00901_ _01155_ VPWR VGND _01293_ sg13g2_o21ai_1
X_07523_ _00863_ _00882_ _01293_ VPWR VGND _01294_ sg13g2_a21oi_1
X_07524_ _01292_ _01294_ _01219_ VPWR VGND _01295_ sg13g2_mux2_1
X_07525_ _00894_ _00861_ VPWR VGND _01296_ sg13g2_nand2_1
X_07526_ _01243_ _01246_ _01003_ _01021_ _01296_ VPWR 
+ VGND
+ _01297_ sg13g2_a221oi_1
X_07527_ _01155_ _00992_ _01215_ _01216_ VPWR VGND 
+ _01298_
+ sg13g2_and4_1
X_07528_ _00861_ _00043_ VPWR VGND _01299_ sg13g2_nor2_1
X_07529_ _00905_ _01209_ _01299_ VPWR VGND _01300_ sg13g2_a21o_1
X_07530_ _01295_ _01297_ _01298_ _01300_ VPWR VGND 
+ _01301_
+ sg13g2_or4_1
X_07531_ _01301_ VPWR VGND _01302_ sg13g2_buf_2
X_07532_ _01288_ _01302_ VPWR VGND _01303_ sg13g2_nor2b_2
X_07533_ _01235_ _01265_ _01026_ VPWR VGND _01304_ sg13g2_o21ai_1
X_07534_ _01303_ _01304_ VPWR VGND _01305_ sg13g2_xnor2_1
X_07535_ _00894_ _01305_ VPWR VGND _01306_ sg13g2_xor2_1
X_07536_ _01282_ _01306_ VPWR VGND _01307_ sg13g2_xnor2_1
X_07537_ _00943_ _01307_ VPWR VGND _01308_ sg13g2_nand2_1
X_07538_ _00093_ _01204_ _01308_ VPWR VGND _01309_ sg13g2_o21ai_1
X_07539_ _01189_ _01309_ VPWR VGND _00145_ sg13g2_nor2_1
X_07540_ _01272_ _01281_ _01305_ VPWR VGND _01310_ sg13g2_o21ai_1
X_07541_ _01272_ _01281_ _01305_ VPWR VGND _01311_ sg13g2_nor3_1
X_07542_ _00894_ _01310_ _01311_ VPWR VGND _01312_ sg13g2_a21oi_1
X_07543_ _00912_ _01153_ VPWR VGND _01313_ sg13g2_nor2_1
X_07544_ _00912_ _01153_ _01284_ _00911_ _01285_ VPWR 
+ VGND
+ _01314_ sg13g2_a221oi_1
X_07545_ _01313_ _01314_ VPWR VGND _01315_ sg13g2_nor2_1
X_07546_ _00915_ \atbs_core_0.adaptive_ctrl_0.n1447_q[3]\ VPWR VGND _01316_ sg13g2_xnor2_1
X_07547_ _01315_ _01316_ VPWR VGND _01317_ sg13g2_xnor2_1
X_07548_ _00923_ \atbs_core_0.adaptive_ctrl_0.spike_i\ _01219_ VPWR VGND _01318_ sg13g2_nor3_1
X_07549_ _01244_ _01246_ _01215_ _01216_ _01006_ VPWR 
+ VGND
+ _01319_ sg13g2_a221oi_1
X_07550_ _01318_ _01319_ _00862_ VPWR VGND _01320_ sg13g2_o21ai_1
X_07551_ _01320_ VPWR VGND _01321_ sg13g2_buf_2
X_07552_ _00992_ _00940_ _00861_ VPWR VGND _01322_ sg13g2_o21ai_1
X_07553_ _01322_ VPWR VGND _01323_ sg13g2_buf_4
X_07554_ _01023_ _01323_ _01161_ VPWR VGND _01324_ sg13g2_o21ai_1
X_07555_ _01324_ VPWR VGND _01325_ sg13g2_buf_2
X_07556_ _01211_ _01321_ _01325_ VPWR VGND _01326_ sg13g2_nand3_1
X_07557_ _01211_ _01317_ _01326_ VPWR VGND _01327_ sg13g2_o21ai_1
X_07558_ _01235_ _01265_ _01303_ VPWR VGND _01328_ sg13g2_nor3_1
X_07559_ _01274_ _01328_ VPWR VGND _01329_ sg13g2_nor2_1
X_07560_ _01327_ _01329_ VPWR VGND _01330_ sg13g2_xnor2_1
X_07561_ _01330_ VPWR VGND _01331_ sg13g2_buf_1
X_07562_ _00893_ _01331_ VPWR VGND _01332_ sg13g2_xnor2_1
X_07563_ _01312_ _01332_ VPWR VGND _01333_ sg13g2_xnor2_1
X_07564_ _00943_ _01333_ VPWR VGND _01334_ sg13g2_nand2_1
X_07565_ _00094_ _01204_ _01334_ VPWR VGND _01335_ sg13g2_o21ai_1
X_07566_ _01189_ _01335_ VPWR VGND _00146_ sg13g2_nor2_1
X_07567_ _01312_ _01331_ _01006_ VPWR VGND _01336_ sg13g2_o21ai_1
X_07568_ _01312_ _01331_ VPWR VGND _01337_ sg13g2_nand2_1
X_07569_ _01336_ _01337_ VPWR VGND _01338_ sg13g2_nand2_1
X_07570_ _00889_ VPWR VGND _01339_ sg13g2_inv_1
X_07571_ _00918_ _01166_ VPWR VGND _01340_ sg13g2_xor2_1
X_07572_ _01313_ _01314_ _01194_ VPWR VGND _01341_ sg13g2_o21ai_1
X_07573_ _01194_ _01313_ _01314_ VPWR VGND _01342_ sg13g2_nor3_1
X_07574_ _00915_ _01341_ _01342_ VPWR VGND _01343_ sg13g2_a21oi_1
X_07575_ _01340_ _01343_ VPWR VGND _01344_ sg13g2_xnor2_1
X_07576_ _01023_ _01323_ VPWR VGND _01345_ sg13g2_nor2_1
X_07577_ _00869_ VPWR VGND _01346_ sg13g2_inv_1
X_07578_ _01346_ \atbs_core_0.adaptive_ctrl_0.spike_i\ _01219_ VPWR VGND _01347_ sg13g2_nor3_1
X_07579_ _01244_ _01246_ _01215_ _01216_ _01339_ VPWR 
+ VGND
+ _01348_ sg13g2_a221oi_1
X_07580_ _01347_ _01348_ _00862_ VPWR VGND _01349_ sg13g2_o21ai_1
X_07581_ _00039_ _01345_ _01349_ VPWR VGND _01350_ sg13g2_o21ai_1
X_07582_ _01350_ VPWR VGND _01351_ sg13g2_buf_1
X_07583_ _01344_ _01351_ _01211_ VPWR VGND _01352_ sg13g2_mux2_1
X_07584_ _01352_ VPWR VGND _01353_ sg13g2_buf_1
X_07585_ _01327_ _01328_ _01274_ VPWR VGND _01354_ sg13g2_a21oi_1
X_07586_ _01353_ _01354_ VPWR VGND _01355_ sg13g2_xnor2_1
X_07587_ _01339_ _01355_ VPWR VGND _01356_ sg13g2_xnor2_1
X_07588_ _01338_ _01356_ VPWR VGND _01357_ sg13g2_xnor2_1
X_07589_ _00943_ _01357_ VPWR VGND _01358_ sg13g2_nand2_1
X_07590_ _00095_ _01204_ _01358_ VPWR VGND _01359_ sg13g2_o21ai_1
X_07591_ _01238_ _01359_ VPWR VGND _00147_ sg13g2_nor2_1
X_07592_ _01355_ VPWR VGND _01360_ sg13g2_inv_1
X_07593_ _01006_ _01331_ _01360_ _01339_ _01312_ VPWR 
+ VGND
+ _01361_ sg13g2_a221oi_1
X_07594_ _01331_ VPWR VGND _01362_ sg13g2_inv_1
X_07595_ _01006_ _01339_ VPWR VGND _01363_ sg13g2_nor2_1
X_07596_ _01006_ _01331_ VPWR VGND _01364_ sg13g2_nor2_1
X_07597_ _00889_ _01355_ VPWR VGND _01365_ sg13g2_and2_1
X_07598_ _01362_ _01363_ _01364_ _01355_ _01365_ VPWR 
+ VGND
+ _01366_ sg13g2_a221oi_1
X_07599_ _01361_ _01366_ VPWR VGND _01367_ sg13g2_nand2b_1
X_07600_ _00868_ VPWR VGND _01368_ sg13g2_inv_1
X_07601_ _01368_ \atbs_core_0.adaptive_ctrl_0.spike_i\ _01219_ VPWR VGND _01369_ sg13g2_nor3_1
X_07602_ _00888_ VPWR VGND _01370_ sg13g2_inv_1
X_07603_ _01244_ _01246_ _01215_ _01216_ _01370_ VPWR 
+ VGND
+ _01371_ sg13g2_a221oi_1
X_07604_ _01369_ _01371_ _00862_ VPWR VGND _01372_ sg13g2_o21ai_1
X_07605_ _00036_ _01345_ _01372_ VPWR VGND _01373_ sg13g2_o21ai_1
X_07606_ _00918_ _01166_ VPWR VGND _01374_ sg13g2_or2_1
X_07607_ _00915_ _01374_ VPWR VGND _01375_ sg13g2_nand2_1
X_07608_ _01375_ VPWR VGND _01376_ sg13g2_inv_1
X_07609_ _00918_ _01166_ VPWR VGND _01377_ sg13g2_and2_1
X_07610_ _01342_ _01374_ _01376_ _01341_ _01377_ VPWR 
+ VGND
+ _01378_ sg13g2_a221oi_1
X_07611_ _00935_ _01173_ VPWR VGND _01379_ sg13g2_xor2_1
X_07612_ _01378_ _01379_ VPWR VGND _01380_ sg13g2_xnor2_1
X_07613_ _01260_ _01380_ VPWR VGND _01381_ sg13g2_and2_1
X_07614_ _01211_ _01373_ _01381_ VPWR VGND _01382_ sg13g2_a21oi_1
X_07615_ _01327_ _01328_ VPWR VGND _01383_ sg13g2_nand2_1
X_07616_ _01353_ _01383_ _01026_ VPWR VGND _01384_ sg13g2_o21ai_1
X_07617_ _01382_ _01384_ VPWR VGND _01385_ sg13g2_xnor2_1
X_07618_ _00888_ _01385_ VPWR VGND _01386_ sg13g2_xnor2_1
X_07619_ _01367_ _01386_ VPWR VGND _01387_ sg13g2_xnor2_1
X_07620_ _00943_ _01387_ VPWR VGND _01388_ sg13g2_nand2_1
X_07621_ _00096_ _01204_ _01388_ VPWR VGND _01389_ sg13g2_o21ai_1
X_07622_ _01238_ _01389_ VPWR VGND _00148_ sg13g2_nor2_1
X_07623_ _00888_ _01385_ VPWR VGND _01390_ sg13g2_or2_1
X_07624_ _00888_ _01385_ VPWR VGND _01391_ sg13g2_nand2_1
X_07625_ _01361_ _01366_ _01391_ VPWR VGND _01392_ sg13g2_nand3b_1
X_07626_ _01390_ _01392_ VPWR VGND _01393_ sg13g2_nand2_1
X_07627_ _00890_ VPWR VGND _01394_ sg13g2_inv_1
X_07628_ _00930_ _01175_ VPWR VGND _01395_ sg13g2_xor2_1
X_07629_ _00935_ _01173_ VPWR VGND _01396_ sg13g2_nor2_1
X_07630_ _00935_ _01173_ VPWR VGND _01397_ sg13g2_nand2_1
X_07631_ _01378_ _01396_ _01397_ VPWR VGND _01398_ sg13g2_o21ai_1
X_07632_ _01395_ _01398_ VPWR VGND _01399_ sg13g2_xnor2_1
X_07633_ _01260_ _01399_ VPWR VGND _01400_ sg13g2_nand2_1
X_07634_ _00873_ _00905_ _00940_ VPWR VGND _01401_ sg13g2_and3_1
X_07635_ _01244_ _01246_ _01215_ _01216_ _01394_ VPWR 
+ VGND
+ _01402_ sg13g2_a221oi_1
X_07636_ _01401_ _01402_ _00862_ VPWR VGND _01403_ sg13g2_o21ai_1
X_07637_ _01023_ _01323_ _01168_ VPWR VGND _01404_ sg13g2_o21ai_1
X_07638_ _01211_ _01403_ _01404_ VPWR VGND _01405_ sg13g2_nand3_1
X_07639_ _01400_ _01405_ VPWR VGND _01406_ sg13g2_and2_1
X_07640_ _01406_ VPWR VGND _01407_ sg13g2_buf_1
X_07641_ _01353_ _01383_ VPWR VGND _01408_ sg13g2_nor2_1
X_07642_ _01382_ _01408_ _01274_ VPWR VGND _01409_ sg13g2_a21oi_1
X_07643_ _01407_ _01409_ VPWR VGND _01410_ sg13g2_xnor2_1
X_07644_ _01394_ _01410_ VPWR VGND _01411_ sg13g2_xnor2_1
X_07645_ _01393_ _01411_ VPWR VGND _01412_ sg13g2_xnor2_1
X_07646_ _00097_ _01204_ _01185_ VPWR VGND _01413_ sg13g2_o21ai_1
X_07647_ _01204_ _01412_ _01413_ VPWR VGND _00149_ sg13g2_a21oi_1
X_07648_ _00943_ _00884_ VPWR VGND _01414_ sg13g2_nand2b_1
X_07649_ _00890_ _01410_ VPWR VGND _01415_ sg13g2_or2_1
X_07650_ _01390_ _01392_ _01415_ VPWR VGND _01416_ sg13g2_nand3_1
X_07651_ _00890_ _01410_ VPWR VGND _01417_ sg13g2_nand2_1
X_07652_ _00926_ \atbs_core_0.adaptive_ctrl_0.n1447_q[7]\ VPWR VGND _01418_ sg13g2_xor2_1
X_07653_ _00930_ _01175_ VPWR VGND _01419_ sg13g2_or2_1
X_07654_ _00930_ _01175_ VPWR VGND _01420_ sg13g2_and2_1
X_07655_ _01398_ _01419_ _01420_ VPWR VGND _01421_ sg13g2_a21oi_1
X_07656_ _01418_ _01421_ VPWR VGND _01422_ sg13g2_xnor2_1
X_07657_ _00034_ \atbs_core_0.adaptive_ctrl_0.spike_i\ _01219_ VPWR VGND _01423_ sg13g2_nor3_1
X_07658_ _01244_ _01246_ _01215_ _01216_ _00033_ VPWR 
+ VGND
+ _01424_ sg13g2_a221oi_1
X_07659_ _01423_ _01424_ _00862_ VPWR VGND _01425_ sg13g2_o21ai_1
X_07660_ _00032_ VPWR VGND _01426_ sg13g2_inv_1
X_07661_ _01023_ _01323_ _01426_ VPWR VGND _01427_ sg13g2_o21ai_1
X_07662_ _01211_ _01425_ _01427_ VPWR VGND _01428_ sg13g2_nand3_1
X_07663_ _01211_ _01422_ _01428_ VPWR VGND _01429_ sg13g2_o21ai_1
X_07664_ _01429_ VPWR VGND _01430_ sg13g2_buf_1
X_07665_ _01026_ _01407_ _01409_ VPWR VGND _01431_ sg13g2_a21oi_1
X_07666_ _01430_ _01431_ VPWR VGND _01432_ sg13g2_xnor2_1
X_07667_ _00033_ _01432_ VPWR VGND _01433_ sg13g2_xor2_1
X_07668_ _01416_ _01417_ _01433_ VPWR VGND _01434_ sg13g2_a21oi_1
X_07669_ _01433_ _01416_ _01417_ VPWR VGND _01435_ sg13g2_nand3_1
X_07670_ _01434_ _01204_ _01435_ VPWR VGND _01436_ sg13g2_nand3b_1
X_07671_ _01414_ _01436_ _01238_ VPWR VGND _00150_ sg13g2_a21oi_1
X_07672_ _00943_ _01185_ VPWR VGND _01437_ sg13g2_nand2_1
X_07673_ _01407_ _01430_ VPWR VGND _01438_ sg13g2_nand2b_1
X_07674_ _01026_ _01438_ _01409_ VPWR VGND _01439_ sg13g2_a21oi_1
X_07675_ _00026_ _01439_ VPWR VGND _01440_ sg13g2_xor2_1
X_07676_ _01437_ _01440_ VPWR VGND _01441_ sg13g2_nor2b_1
X_07677_ _01434_ _01441_ VPWR VGND _01442_ sg13g2_nand2_1
X_07678_ _00884_ _01432_ VPWR VGND _01443_ sg13g2_and2_1
X_07679_ _01434_ _01437_ _01440_ _01443_ VPWR VGND 
+ _01444_
+ sg13g2_or4_1
X_07680_ _01443_ _01441_ VPWR VGND _01445_ sg13g2_nand2_1
X_07681_ _00943_ _01185_ _00885_ VPWR VGND _01446_ sg13g2_nand3b_1
X_07682_ _01442_ _01444_ _01445_ _01446_ VPWR VGND 
+ _00151_
+ sg13g2_nand4_1
X_07683_ _01029_ VPWR VGND _01447_ sg13g2_buf_1
X_07684_ _00992_ _01003_ _01021_ _01206_ VPWR VGND 
+ _01448_
+ sg13g2_nand4_1
X_07685_ _01448_ VPWR VGND _01449_ sg13g2_buf_2
X_07686_ _01109_ _01449_ _00862_ VPWR VGND _01450_ sg13g2_o21ai_1
X_07687_ _01230_ _01449_ VPWR VGND _01451_ sg13g2_nor2_1
X_07688_ _01224_ _01449_ _01450_ _01212_ _01451_ VPWR 
+ VGND
+ _01452_ sg13g2_a221oi_1
X_07689_ _01452_ VPWR VGND _01453_ sg13g2_buf_4
X_07690_ _00909_ _01453_ VPWR VGND _01454_ sg13g2_xnor2_1
X_07691_ _01447_ _01454_ VPWR VGND _01455_ sg13g2_nor2_1
X_07692_ _00098_ _01447_ _01455_ VPWR VGND _01456_ sg13g2_a21oi_1
X_07693_ _01238_ _01456_ VPWR VGND _00152_ sg13g2_nor2_1
X_07694_ _00860_ \atbs_core_0.adaptive_ctrl_0.spike_i\ VPWR VGND _01457_ sg13g2_nor2_1
X_07695_ _01457_ VPWR VGND _01458_ sg13g2_buf_2
X_07696_ _00909_ _01458_ VPWR VGND _01459_ sg13g2_xnor2_1
X_07697_ _01453_ _01459_ VPWR VGND _01460_ sg13g2_nand2_1
X_07698_ _00992_ _01215_ _01216_ _01206_ VPWR VGND 
+ _01461_
+ sg13g2_and4_1
X_07699_ _01461_ VPWR VGND _01462_ sg13g2_buf_4
X_07700_ _00907_ _00860_ \atbs_core_0.adaptive_ctrl_0.spike_i\ _01219_ VPWR VGND 
+ _01463_
+ sg13g2_nor4_2
X_07701_ _00861_ _01241_ VPWR VGND _01464_ sg13g2_nand2_1
X_07702_ _01244_ _01246_ _01215_ _01216_ _01464_ VPWR 
+ VGND
+ _01465_ sg13g2_a221oi_1
X_07703_ _01462_ _01463_ _01465_ VPWR VGND _01466_ sg13g2_nor3_1
X_07704_ _01023_ _01323_ _01148_ VPWR VGND _01467_ sg13g2_o21ai_1
X_07705_ _01467_ VPWR VGND _01468_ sg13g2_buf_4
X_07706_ _01262_ _01462_ _01466_ _01468_ VPWR VGND 
+ _01469_
+ sg13g2_a22oi_1
X_07707_ _01469_ VPWR VGND _01470_ sg13g2_buf_2
X_07708_ _00907_ _01470_ VPWR VGND _01471_ sg13g2_xnor2_1
X_07709_ _01460_ _01471_ VPWR VGND _01472_ sg13g2_xnor2_1
X_07710_ _01447_ _01472_ VPWR VGND _01473_ sg13g2_nor2_1
X_07711_ _00099_ _01447_ _01473_ VPWR VGND _01474_ sg13g2_a21oi_1
X_07712_ _01238_ _01474_ VPWR VGND _00153_ sg13g2_nor2_1
X_07713_ _01262_ _01462_ _01466_ _01468_ _01458_ VPWR 
+ VGND
+ _01475_ sg13g2_a221oi_1
X_07714_ _01458_ _01466_ _01468_ VPWR VGND _01476_ sg13g2_and3_1
X_07715_ _01475_ _01476_ _00872_ VPWR VGND _01477_ sg13g2_o21ai_1
X_07716_ _00872_ _01476_ _00871_ VPWR VGND _01478_ sg13g2_o21ai_1
X_07717_ _01453_ VPWR VGND _01479_ sg13g2_inv_1
X_07718_ _01477_ _01478_ _01479_ VPWR VGND _01480_ sg13g2_a21o_1
X_07719_ _01458_ _01453_ VPWR VGND _01481_ sg13g2_nand2_1
X_07720_ _00871_ _01470_ _01481_ VPWR VGND _01482_ sg13g2_nand3_1
X_07721_ _01480_ _01482_ VPWR VGND _01483_ sg13g2_nand2_1
X_07722_ _01295_ _01297_ _01298_ _01299_ VPWR VGND 
+ _01484_
+ sg13g2_nor4_1
X_07723_ _01287_ _01449_ VPWR VGND _01485_ sg13g2_nor2_1
X_07724_ _01484_ _01449_ _01485_ VPWR VGND _01486_ sg13g2_a21oi_1
X_07725_ _01486_ VPWR VGND _01487_ sg13g2_buf_4
X_07726_ _01453_ _01470_ _01458_ VPWR VGND _01488_ sg13g2_o21ai_1
X_07727_ _01487_ _01488_ VPWR VGND _01489_ sg13g2_xnor2_1
X_07728_ _00877_ _01489_ VPWR VGND _01490_ sg13g2_xnor2_1
X_07729_ _01483_ _01490_ VPWR VGND _01491_ sg13g2_xnor2_1
X_07730_ _01447_ _01491_ VPWR VGND _01492_ sg13g2_nor2_1
X_07731_ _00100_ _01447_ _01492_ VPWR VGND _01493_ sg13g2_a21oi_1
X_07732_ _01238_ _01493_ VPWR VGND _00154_ sg13g2_nor2_1
X_07733_ _01289_ _01480_ _01482_ VPWR VGND _01494_ sg13g2_nand3_1
X_07734_ _01480_ _01482_ _01289_ VPWR VGND _01495_ sg13g2_a21oi_1
X_07735_ _01489_ _01494_ _01495_ VPWR VGND _01496_ sg13g2_a21o_1
X_07736_ _01321_ _01325_ VPWR VGND _01497_ sg13g2_nand2_1
X_07737_ _01449_ VPWR VGND _01498_ sg13g2_buf_2
X_07738_ _01317_ _01497_ _01498_ VPWR VGND _01499_ sg13g2_mux2_1
X_07739_ _01499_ VPWR VGND _01500_ sg13g2_buf_1
X_07740_ _01453_ _01470_ _01487_ VPWR VGND _01501_ sg13g2_or3_1
X_07741_ _01501_ VPWR VGND _01502_ sg13g2_buf_2
X_07742_ _01458_ _01502_ VPWR VGND _01503_ sg13g2_nand2_1
X_07743_ _01500_ _01503_ VPWR VGND _01504_ sg13g2_xnor2_1
X_07744_ _00876_ _01504_ VPWR VGND _01505_ sg13g2_xnor2_1
X_07745_ _01496_ _01505_ VPWR VGND _01506_ sg13g2_xnor2_1
X_07746_ _01029_ _01506_ VPWR VGND _01507_ sg13g2_nor2_1
X_07747_ _00101_ _01447_ _01507_ VPWR VGND _01508_ sg13g2_a21oi_1
X_07748_ _01238_ _01508_ VPWR VGND _00155_ sg13g2_nor2_1
X_07749_ _00876_ _01504_ VPWR VGND _01509_ sg13g2_nor2_1
X_07750_ _01489_ _01494_ _01504_ _00876_ _01495_ VPWR 
+ VGND
+ _01510_ sg13g2_a221oi_1
X_07751_ _01510_ VPWR VGND _01511_ sg13g2_buf_1
X_07752_ _01509_ _01511_ VPWR VGND _01512_ sg13g2_nor2_2
X_07753_ _01344_ _01351_ _01498_ VPWR VGND _01513_ sg13g2_mux2_1
X_07754_ _01513_ VPWR VGND _01514_ sg13g2_buf_1
X_07755_ _01500_ _01502_ _01458_ VPWR VGND _01515_ sg13g2_o21ai_1
X_07756_ _01514_ _01515_ VPWR VGND _01516_ sg13g2_xor2_1
X_07757_ _01346_ _01516_ VPWR VGND _01517_ sg13g2_xnor2_1
X_07758_ _01512_ _01517_ VPWR VGND _01518_ sg13g2_xnor2_1
X_07759_ _01029_ _01518_ VPWR VGND _01519_ sg13g2_nor2_1
X_07760_ _00102_ _01447_ _01519_ VPWR VGND _01520_ sg13g2_a21oi_1
X_07761_ _01238_ _01520_ VPWR VGND _00156_ sg13g2_nor2_1
X_07762_ _01509_ _01511_ _01516_ VPWR VGND _01521_ sg13g2_nor3_2
X_07763_ _01509_ _01511_ _01516_ VPWR VGND _01522_ sg13g2_o21ai_1
X_07764_ _00869_ _01521_ _01522_ VPWR VGND _01523_ sg13g2_o21ai_1
X_07765_ _01380_ _01373_ _01498_ VPWR VGND _01524_ sg13g2_mux2_1
X_07766_ _01500_ _01502_ _01514_ VPWR VGND _01525_ sg13g2_nor3_1
X_07767_ _00906_ _01525_ VPWR VGND _01526_ sg13g2_nor2_1
X_07768_ _01524_ _01526_ VPWR VGND _01527_ sg13g2_xnor2_1
X_07769_ _01527_ VPWR VGND _01528_ sg13g2_buf_1
X_07770_ _00868_ _01528_ VPWR VGND _01529_ sg13g2_xnor2_1
X_07771_ _01523_ _01529_ VPWR VGND _01530_ sg13g2_xnor2_1
X_07772_ _00103_ _01029_ VPWR VGND _01531_ sg13g2_nand2_1
X_07773_ _01447_ _01530_ _01531_ VPWR VGND _01532_ sg13g2_o21ai_1
X_07774_ _01185_ _01532_ VPWR VGND _00157_ sg13g2_and2_1
X_07775_ _00104_ _01447_ VPWR VGND _01533_ sg13g2_nand2_1
X_07776_ _01523_ _01528_ _01368_ VPWR VGND _01534_ sg13g2_o21ai_1
X_07777_ _01523_ _01528_ VPWR VGND _01535_ sg13g2_nand2_1
X_07778_ _01399_ _01462_ VPWR VGND _01536_ sg13g2_nand2_1
X_07779_ _01403_ _01404_ _01498_ VPWR VGND _01537_ sg13g2_nand3_1
X_07780_ _01536_ _01537_ VPWR VGND _01538_ sg13g2_and2_1
X_07781_ _01538_ VPWR VGND _01539_ sg13g2_buf_1
X_07782_ _01500_ _01502_ _01514_ _01524_ VPWR VGND 
+ _01540_
+ sg13g2_nor4_1
X_07783_ _00906_ _01540_ VPWR VGND _01541_ sg13g2_nor2_1
X_07784_ _01539_ _01541_ VPWR VGND _01542_ sg13g2_xor2_1
X_07785_ _00873_ _01542_ VPWR VGND _01543_ sg13g2_nand2_1
X_07786_ _01543_ VPWR VGND _01544_ sg13g2_inv_1
X_07787_ _00873_ _01542_ VPWR VGND _01545_ sg13g2_nor2_1
X_07788_ _01544_ _01545_ VPWR VGND _01546_ sg13g2_nor2_1
X_07789_ _01534_ _01535_ _01546_ VPWR VGND _01547_ sg13g2_a21oi_1
X_07790_ _01546_ _01534_ _01535_ VPWR VGND _01548_ sg13g2_and3_1
X_07791_ _01547_ _01548_ _01030_ VPWR VGND _01549_ sg13g2_o21ai_1
X_07792_ _01533_ _01549_ _01238_ VPWR VGND _00158_ sg13g2_a21oi_1
X_07793_ _01540_ VPWR VGND _01550_ sg13g2_inv_1
X_07794_ _01539_ _01550_ _01458_ VPWR VGND _01551_ sg13g2_o21ai_1
X_07795_ _01551_ VPWR VGND _01552_ sg13g2_buf_1
X_07796_ _01425_ _01427_ _01498_ VPWR VGND _01553_ sg13g2_nand3_1
X_07797_ _01422_ _01498_ _01553_ VPWR VGND _01554_ sg13g2_o21ai_1
X_07798_ _01554_ VPWR VGND _01555_ sg13g2_buf_1
X_07799_ _01552_ _01555_ VPWR VGND _01556_ sg13g2_xor2_1
X_07800_ _00925_ _01095_ VPWR VGND _01557_ sg13g2_nor2_1
X_07801_ _01556_ _01557_ VPWR VGND _01558_ sg13g2_nand2_1
X_07802_ _00878_ _01029_ _01095_ VPWR VGND _01559_ sg13g2_nor3_1
X_07803_ _01543_ _01556_ _01559_ VPWR VGND _01560_ sg13g2_nand3_1
X_07804_ _00869_ _01512_ VPWR VGND _01561_ sg13g2_nor2_1
X_07805_ _01528_ _01561_ _01368_ VPWR VGND _01562_ sg13g2_o21ai_1
X_07806_ _00869_ _01521_ VPWR VGND _01563_ sg13g2_nor2_1
X_07807_ _01368_ _01528_ VPWR VGND _01564_ sg13g2_nor2_1
X_07808_ _01512_ _01564_ _00870_ VPWR VGND _01565_ sg13g2_o21ai_1
X_07809_ _01563_ _01528_ _01565_ _01516_ _01545_ VPWR 
+ VGND
+ _01566_ sg13g2_a221oi_1
X_07810_ _01562_ _01566_ VPWR VGND _01567_ sg13g2_nand2_1
X_07811_ _01558_ _01560_ _01567_ VPWR VGND _01568_ sg13g2_mux2_1
X_07812_ _01552_ _01555_ VPWR VGND _01569_ sg13g2_xnor2_1
X_07813_ _01543_ _01569_ _01567_ _01557_ VPWR VGND 
+ _01570_
+ sg13g2_nand4_1
X_07814_ _01569_ _01562_ _01566_ _01559_ VPWR VGND 
+ _01571_
+ sg13g2_nand4_1
X_07815_ _01543_ _01556_ VPWR VGND _01572_ sg13g2_nor2_1
X_07816_ _00925_ _01095_ _01543_ _01569_ VPWR VGND 
+ _01573_
+ sg13g2_nor4_1
X_07817_ _01029_ _01557_ _01572_ _01559_ _01573_ VPWR 
+ VGND
+ _01574_ sg13g2_a221oi_1
X_07818_ _01568_ _01570_ _01571_ _01574_ VPWR VGND 
+ _00159_
+ sg13g2_nand4_1
X_07819_ _01562_ _01566_ _01544_ VPWR VGND _01575_ sg13g2_a21oi_1
X_07820_ _01552_ _01555_ VPWR VGND _01576_ sg13g2_nand2_1
X_07821_ _01458_ _01552_ _01555_ VPWR VGND _01577_ sg13g2_a21o_1
X_07822_ _00034_ _01577_ VPWR VGND _01578_ sg13g2_nand2b_1
X_07823_ _00034_ _00906_ VPWR VGND _01579_ sg13g2_nand2_1
X_07824_ _01030_ _01576_ _01578_ _01579_ VPWR VGND 
+ _01580_
+ sg13g2_nand4_1
X_07825_ _00874_ _01185_ _01575_ _01580_ VPWR VGND 
+ _01581_
+ sg13g2_nand4_1
X_07826_ _00874_ _01095_ _01580_ VPWR VGND _01582_ sg13g2_nor3_1
X_07827_ _01575_ _01582_ VPWR VGND _01583_ sg13g2_nand2_1
X_07828_ _00878_ _01577_ VPWR VGND _01584_ sg13g2_nor2_1
X_07829_ _00862_ _00905_ _01553_ VPWR VGND _01585_ sg13g2_nand3_1
X_07830_ _01552_ _01585_ _00034_ VPWR VGND _01586_ sg13g2_a21oi_1
X_07831_ _01552_ _01579_ _01555_ VPWR VGND _01587_ sg13g2_a21oi_1
X_07832_ _00925_ _01586_ _01587_ VPWR VGND _01588_ sg13g2_nor3_1
X_07833_ _01584_ _01588_ _01030_ VPWR VGND _01589_ sg13g2_o21ai_1
X_07834_ _00874_ _01185_ _01589_ VPWR VGND _01590_ sg13g2_nand3_1
X_07835_ _01589_ _01185_ _00927_ VPWR VGND _01591_ sg13g2_nand3b_1
X_07836_ _01590_ _01591_ _01575_ VPWR VGND _01592_ sg13g2_a21o_1
X_07837_ _01581_ _01583_ _01592_ VPWR VGND _00160_ sg13g2_nand3_1
X_07838_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[16]\ VPWR VGND _01593_ sg13g2_buf_1
X_07839_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[15]\ VPWR VGND _01594_ sg13g2_buf_1
X_07840_ _01594_ VPWR VGND _01595_ sg13g2_buf_1
X_07841_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[15]\ VPWR VGND _01596_ sg13g2_buf_1
X_07842_ _01595_ _01596_ VPWR VGND _01597_ sg13g2_nor2_1
X_07843_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[14]\ VPWR VGND _01598_ sg13g2_buf_1
X_07844_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[13]\ VPWR VGND _01599_ sg13g2_buf_1
X_07845_ _01599_ VPWR VGND _01600_ sg13g2_inv_1
X_07846_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[10]\ VPWR VGND _01601_ sg13g2_buf_1
X_07847_ _01601_ VPWR VGND _01602_ sg13g2_inv_1
X_07848_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[9]\ VPWR VGND _01603_ sg13g2_buf_1
X_07849_ _01603_ VPWR VGND _01604_ sg13g2_buf_2
X_07850_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[8]\ VPWR VGND _01605_ sg13g2_buf_1
X_07851_ _01605_ VPWR VGND _01606_ sg13g2_buf_2
X_07852_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[8]\ VPWR VGND _01607_ sg13g2_buf_1
X_07853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[6]\ VPWR VGND _01608_ sg13g2_buf_4
X_07854_ _01608_ VPWR VGND _01609_ sg13g2_buf_4
X_07855_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[6]\ VPWR VGND _01610_ sg13g2_buf_1
X_07856_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[7]\ VPWR VGND _01611_ sg13g2_buf_1
X_07857_ _01609_ _01610_ _01611_ VPWR VGND _01612_ sg13g2_a21o_1
X_07858_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[7]\ VPWR VGND _01613_ sg13g2_buf_2
X_07859_ _01613_ VPWR VGND _01614_ sg13g2_buf_2
X_07860_ _01609_ _01611_ _01610_ VPWR VGND _01615_ sg13g2_and3_1
X_07861_ _01615_ VPWR VGND _01616_ sg13g2_buf_1
X_07862_ _01606_ _01607_ _01612_ _01614_ _01616_ VPWR 
+ VGND
+ _01617_ sg13g2_a221oi_1
X_07863_ _01617_ VPWR VGND _01618_ sg13g2_buf_1
X_07864_ _01606_ VPWR VGND _01619_ sg13g2_buf_2
X_07865_ _01619_ _01607_ VPWR VGND _01620_ sg13g2_nor2_1
X_07866_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[9]\ VPWR VGND _01621_ sg13g2_buf_1
X_07867_ _01621_ VPWR VGND _01622_ sg13g2_inv_1
X_07868_ _01618_ _01620_ _01622_ VPWR VGND _01623_ sg13g2_o21ai_1
X_07869_ _01623_ VPWR VGND _01624_ sg13g2_buf_1
X_07870_ _01622_ _01618_ _01620_ VPWR VGND _01625_ sg13g2_nor3_1
X_07871_ _01604_ _01624_ _01625_ VPWR VGND _01626_ sg13g2_a21oi_1
X_07872_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[10]\ VPWR VGND _01627_ sg13g2_buf_1
X_07873_ _01627_ VPWR VGND _01628_ sg13g2_inv_1
X_07874_ _01602_ _01626_ _01628_ VPWR VGND _01629_ sg13g2_o21ai_1
X_07875_ _01629_ VPWR VGND _01630_ sg13g2_buf_2
X_07876_ _01602_ _01626_ VPWR VGND _01631_ sg13g2_nand2_1
X_07877_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[13]\ VPWR VGND _01632_ sg13g2_buf_1
X_07878_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[11]\ VPWR VGND _01633_ sg13g2_buf_1
X_07879_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[12]\ VPWR VGND _01634_ sg13g2_buf_1
X_07880_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[12]\ VPWR VGND _01635_ sg13g2_buf_1
X_07881_ _01634_ _01635_ VPWR VGND _01636_ sg13g2_and2_1
X_07882_ _01636_ VPWR VGND _01637_ sg13g2_buf_1
X_07883_ _01632_ _01633_ _01637_ VPWR VGND _01638_ sg13g2_or3_1
X_07884_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[11]\ VPWR VGND _01639_ sg13g2_buf_1
X_07885_ _01639_ _01632_ _01637_ VPWR VGND _01640_ sg13g2_or3_1
X_07886_ _01630_ _01631_ _01638_ _01640_ VPWR VGND 
+ _01641_
+ sg13g2_a22oi_1
X_07887_ _01634_ _01635_ VPWR VGND _01642_ sg13g2_or2_1
X_07888_ _01642_ VPWR VGND _01643_ sg13g2_buf_1
X_07889_ _01632_ _01643_ VPWR VGND _01644_ sg13g2_nor2_1
X_07890_ _01633_ _01640_ VPWR VGND _01645_ sg13g2_nor2_1
X_07891_ _01600_ _01641_ _01644_ _01645_ VPWR VGND 
+ _01646_
+ sg13g2_nor4_2
X_07892_ _01604_ _01624_ _01625_ VPWR VGND _01647_ sg13g2_a21o_1
X_07893_ _01627_ VPWR VGND _01648_ sg13g2_buf_1
X_07894_ _01601_ _01647_ _01648_ VPWR VGND _01649_ sg13g2_a21oi_1
X_07895_ _01601_ _01647_ VPWR VGND _01650_ sg13g2_nor2_1
X_07896_ _01632_ _01633_ _01643_ VPWR VGND _01651_ sg13g2_nand3_1
X_07897_ _01649_ _01650_ _01651_ VPWR VGND _01652_ sg13g2_nor3_1
X_07898_ _01639_ _01632_ _01643_ VPWR VGND _01653_ sg13g2_and3_1
X_07899_ _01630_ _01631_ _01653_ VPWR VGND _01654_ sg13g2_nand3_1
X_07900_ _01632_ _01637_ _01653_ _01633_ VPWR VGND 
+ _01655_
+ sg13g2_a22oi_1
X_07901_ _01652_ _01654_ _01655_ VPWR VGND _01656_ sg13g2_nand3b_1
X_07902_ _01596_ _01598_ _01646_ _01656_ VPWR VGND 
+ _01657_
+ sg13g2_nor4_1
X_07903_ _01594_ VPWR VGND _01658_ sg13g2_buf_1
X_07904_ _01658_ _01598_ _01646_ _01656_ VPWR VGND 
+ _01659_
+ sg13g2_nor4_1
X_07905_ _01657_ _01659_ VPWR VGND _01660_ sg13g2_or2_1
X_07906_ _01634_ VPWR VGND _01661_ sg13g2_buf_1
X_07907_ _01661_ VPWR VGND _01662_ sg13g2_buf_1
X_07908_ _01662_ _01635_ VPWR VGND _01663_ sg13g2_nor2_1
X_07909_ _01633_ VPWR VGND _01664_ sg13g2_inv_1
X_07910_ _01649_ _01650_ _01664_ VPWR VGND _01665_ sg13g2_o21ai_1
X_07911_ _01639_ VPWR VGND _01666_ sg13g2_buf_1
X_07912_ _01666_ VPWR VGND _01667_ sg13g2_buf_1
X_07913_ _01664_ _01649_ _01650_ VPWR VGND _01668_ sg13g2_nor3_1
X_07914_ _01662_ _01635_ _01665_ _01667_ _01668_ VPWR 
+ VGND
+ _01669_ sg13g2_a221oi_1
X_07915_ _01663_ _01669_ VPWR VGND _01670_ sg13g2_nor2_1
X_07916_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[14]\ VPWR VGND _01671_ sg13g2_buf_1
X_07917_ _01671_ VPWR VGND _01672_ sg13g2_buf_1
X_07918_ _01672_ _01596_ VPWR VGND _01673_ sg13g2_or2_1
X_07919_ _01658_ VPWR VGND _01674_ sg13g2_inv_1
X_07920_ _01672_ VPWR VGND _01675_ sg13g2_inv_1
X_07921_ _01674_ _01675_ VPWR VGND _01676_ sg13g2_nand2_1
X_07922_ _01632_ _01670_ _01673_ _01676_ _01646_ VPWR 
+ VGND
+ _01677_ sg13g2_a221oi_1
X_07923_ _01673_ _01676_ _01598_ VPWR VGND _01678_ sg13g2_a21oi_1
X_07924_ _01597_ _01660_ _01677_ _01678_ VPWR VGND 
+ _01679_
+ sg13g2_nor4_2
X_07925_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[16]\ VPWR VGND _01680_ sg13g2_buf_1
X_07926_ _01680_ VPWR VGND _01681_ sg13g2_buf_1
X_07927_ _01681_ VPWR VGND _01682_ sg13g2_buf_1
X_07928_ _01593_ _01679_ _01682_ VPWR VGND _01683_ sg13g2_a21o_1
X_07929_ _01593_ _01679_ _01683_ VPWR VGND _01684_ sg13g2_o21ai_1
X_07930_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[17]\ VPWR VGND _01685_ sg13g2_buf_1
X_07931_ _01685_ VPWR VGND _01686_ sg13g2_buf_1
X_07932_ _01686_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[17]\ VPWR VGND _01687_ sg13g2_xor2_1
X_07933_ _01684_ _01687_ VPWR VGND _01688_ sg13g2_xnor2_1
X_07934_ _00020_ VPWR VGND _01689_ sg13g2_buf_1
X_07935_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[17]\ VPWR VGND _01690_ sg13g2_buf_1
X_07936_ _01689_ _01690_ VPWR VGND _01691_ sg13g2_nor2_1
X_07937_ _01691_ VPWR VGND _01692_ sg13g2_inv_1
X_07938_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2072_o\ VPWR VGND _01693_ sg13g2_inv_1
X_07939_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[17]\ VPWR VGND _01694_ sg13g2_inv_1
X_07940_ _01694_ _01684_ VPWR VGND _01695_ sg13g2_nor2_1
X_07941_ _01685_ VPWR VGND _01696_ sg13g2_inv_1
X_07942_ _01696_ VPWR VGND _01697_ sg13g2_buf_1
X_07943_ _01697_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2072_o\ VPWR VGND _01698_ sg13g2_nor2_1
X_07944_ _01694_ _01684_ VPWR VGND _01699_ sg13g2_nand2_1
X_07945_ _01693_ _01695_ _01698_ _01699_ VPWR VGND 
+ _01700_
+ sg13g2_a22oi_1
X_07946_ _01688_ _01692_ _01700_ VPWR VGND _01701_ sg13g2_o21ai_1
X_07947_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[14]\ VPWR VGND _01702_ sg13g2_buf_1
X_07948_ _01702_ VPWR VGND _01703_ sg13g2_inv_1
X_07949_ _01646_ _01656_ VPWR VGND _01704_ sg13g2_or2_1
X_07950_ _01704_ VPWR VGND _01705_ sg13g2_buf_1
X_07951_ _01672_ VPWR VGND _01706_ sg13g2_buf_1
X_07952_ _01706_ _01598_ VPWR VGND _01707_ sg13g2_xnor2_1
X_07953_ _01705_ _01707_ VPWR VGND _01708_ sg13g2_xnor2_1
X_07954_ _00013_ VPWR VGND _01709_ sg13g2_buf_1
X_07955_ _01709_ _01708_ VPWR VGND _01710_ sg13g2_xnor2_1
X_07956_ _01599_ VPWR VGND _01711_ sg13g2_buf_1
X_07957_ _01711_ VPWR VGND _01712_ sg13g2_buf_1
X_07958_ _01712_ VPWR VGND _01713_ sg13g2_buf_1
X_07959_ _01713_ _01632_ VPWR VGND _01714_ sg13g2_xor2_1
X_07960_ _01663_ _01669_ _01714_ VPWR VGND _01715_ sg13g2_or3_1
X_07961_ _01663_ _01669_ _01714_ VPWR VGND _01716_ sg13g2_o21ai_1
X_07962_ _01667_ VPWR VGND _01717_ sg13g2_buf_1
X_07963_ _01717_ _01665_ _01668_ VPWR VGND _01718_ sg13g2_a21oi_1
X_07964_ _01662_ VPWR VGND _01719_ sg13g2_buf_1
X_07965_ _01719_ _01635_ VPWR VGND _01720_ sg13g2_xnor2_1
X_07966_ _01718_ _01720_ VPWR VGND _01721_ sg13g2_xnor2_1
X_07967_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[12]\ VPWR VGND _01722_ sg13g2_buf_1
X_07968_ _01715_ _01716_ _01721_ _01722_ VPWR VGND 
+ _01723_
+ sg13g2_a22oi_1
X_07969_ _00014_ VPWR VGND _01724_ sg13g2_buf_1
X_07970_ _01724_ VPWR VGND _01725_ sg13g2_inv_1
X_07971_ _01722_ _01721_ _01725_ VPWR VGND _01726_ sg13g2_a21oi_1
X_07972_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[10]\ VPWR VGND _01727_ sg13g2_buf_1
X_07973_ _01727_ VPWR VGND _01728_ sg13g2_inv_1
X_07974_ _01648_ VPWR VGND _01729_ sg13g2_buf_1
X_07975_ _01729_ VPWR VGND _01730_ sg13g2_buf_1
X_07976_ _01730_ _01601_ VPWR VGND _01731_ sg13g2_xor2_1
X_07977_ _01626_ _01731_ VPWR VGND _01732_ sg13g2_xnor2_1
X_07978_ _01728_ _01732_ VPWR VGND _01733_ sg13g2_nor2_1
X_07979_ _01618_ _01620_ VPWR VGND _01734_ sg13g2_nor2_1
X_07980_ _01604_ VPWR VGND _01735_ sg13g2_buf_1
X_07981_ _01735_ VPWR VGND _01736_ sg13g2_buf_1
X_07982_ _01736_ _01621_ VPWR VGND _01737_ sg13g2_xor2_1
X_07983_ _00018_ VPWR VGND _01738_ sg13g2_buf_1
X_07984_ _01738_ VPWR VGND _01739_ sg13g2_buf_1
X_07985_ _01736_ VPWR VGND _01740_ sg13g2_buf_1
X_07986_ _01740_ _01621_ VPWR VGND _01741_ sg13g2_nand2_1
X_07987_ _01739_ _01734_ _01741_ VPWR VGND _01742_ sg13g2_a21oi_1
X_07988_ _01734_ _01737_ _01742_ VPWR VGND _01743_ sg13g2_a21oi_1
X_07989_ _01603_ VPWR VGND _01744_ sg13g2_inv_1
X_07990_ _01739_ _01625_ _01624_ VPWR VGND _01745_ sg13g2_o21ai_1
X_07991_ _01739_ _01624_ VPWR VGND _01746_ sg13g2_nor2_1
X_07992_ _01744_ _01745_ _01746_ VPWR VGND _01747_ sg13g2_a21oi_1
X_07993_ _00017_ VPWR VGND _01748_ sg13g2_buf_1
X_07994_ _01627_ _01748_ VPWR VGND _01749_ sg13g2_xnor2_1
X_07995_ _01749_ VPWR VGND _01750_ sg13g2_buf_1
X_07996_ _01601_ _01750_ VPWR VGND _01751_ sg13g2_xnor2_1
X_07997_ _01743_ _01747_ _01751_ VPWR VGND _01752_ sg13g2_mux2_1
X_07998_ _01619_ VPWR VGND _01753_ sg13g2_buf_2
X_07999_ _00019_ VPWR VGND _01754_ sg13g2_buf_1
X_08000_ _01753_ _01754_ VPWR VGND _01755_ sg13g2_xnor2_1
X_08001_ _01755_ VPWR VGND _01756_ sg13g2_buf_2
X_08002_ _01607_ _01756_ VPWR VGND _01757_ sg13g2_xor2_1
X_08003_ _01614_ VPWR VGND _01758_ sg13g2_buf_1
X_08004_ _01758_ VPWR VGND _01759_ sg13g2_buf_1
X_08005_ _00010_ VPWR VGND _01760_ sg13g2_buf_1
X_08006_ _01760_ VPWR VGND _01761_ sg13g2_buf_1
X_08007_ _01611_ VPWR VGND _01762_ sg13g2_buf_1
X_08008_ _01608_ VPWR VGND _01763_ sg13g2_buf_2
X_08009_ _01763_ VPWR VGND _01764_ sg13g2_buf_2
X_08010_ _01764_ _01610_ VPWR VGND _01765_ sg13g2_nand2_1
X_08011_ _01761_ _01762_ _01765_ VPWR VGND _01766_ sg13g2_a21oi_1
X_08012_ _01758_ VPWR VGND _01767_ sg13g2_buf_1
X_08013_ _01767_ _01765_ VPWR VGND _01768_ sg13g2_xnor2_1
X_08014_ _01759_ _01766_ _01768_ _01762_ VPWR VGND 
+ _01769_
+ sg13g2_a22oi_1
X_08015_ _01610_ VPWR VGND _01770_ sg13g2_buf_1
X_08016_ _00011_ VPWR VGND _01771_ sg13g2_buf_1
X_08017_ _01764_ _01771_ VPWR VGND _01772_ sg13g2_xnor2_1
X_08018_ _01772_ VPWR VGND _01773_ sg13g2_buf_1
X_08019_ _01773_ VPWR VGND _01774_ sg13g2_buf_1
X_08020_ _01770_ _01774_ VPWR VGND _01775_ sg13g2_or2_1
X_08021_ _01770_ _01774_ VPWR VGND _01776_ sg13g2_nand2_1
X_08022_ _01761_ _01762_ VPWR VGND _01777_ sg13g2_nor2_1
X_08023_ _01761_ _01616_ _01612_ VPWR VGND _01778_ sg13g2_o21ai_1
X_08024_ _01613_ VPWR VGND _01779_ sg13g2_inv_1
X_08025_ _01779_ VPWR VGND _01780_ sg13g2_buf_2
X_08026_ _01765_ _01777_ _01778_ _01780_ _01757_ VPWR 
+ VGND
+ _01781_ sg13g2_a221oi_1
X_08027_ _01757_ _01769_ _01775_ _01776_ _01781_ VPWR 
+ VGND
+ _01782_ sg13g2_a221oi_1
X_08028_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[4]\ VPWR VGND _01783_ sg13g2_buf_1
X_08029_ _01783_ VPWR VGND _01784_ sg13g2_buf_1
X_08030_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[4]\ VPWR VGND _01785_ sg13g2_inv_1
X_08031_ _01784_ _01785_ VPWR VGND _01786_ sg13g2_nor2_1
X_08032_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[2]\ VPWR VGND _01787_ sg13g2_buf_1
X_08033_ _01787_ VPWR VGND _01788_ sg13g2_buf_1
X_08034_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[2]\ VPWR VGND _01789_ sg13g2_inv_1
X_08035_ _01788_ _01789_ VPWR VGND _01790_ sg13g2_nor2_1
X_08036_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[0]\ VPWR VGND _01791_ sg13g2_buf_1
X_08037_ _01791_ VPWR VGND _01792_ sg13g2_buf_1
X_08038_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ VPWR VGND _01793_ sg13g2_nor2b_1
X_08039_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _01793_ VPWR VGND _01794_ sg13g2_nand2_1
X_08040_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[1]\ VPWR VGND _01795_ sg13g2_buf_1
X_08041_ _01795_ VPWR VGND _01796_ sg13g2_inv_1
X_08042_ _01796_ VPWR VGND _01797_ sg13g2_buf_1
X_08043_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _01793_ _01797_ VPWR VGND _01798_ sg13g2_o21ai_1
X_08044_ _01788_ _01789_ _01794_ _01798_ VPWR VGND 
+ _01799_
+ sg13g2_a22oi_1
X_08045_ _01790_ _01799_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ VPWR VGND _01800_ sg13g2_o21ai_1
X_08046_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[3]\ VPWR VGND _01801_ sg13g2_buf_1
X_08047_ _01801_ VPWR VGND _01802_ sg13g2_buf_1
X_08048_ _01802_ VPWR VGND _01803_ sg13g2_buf_1
X_08049_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _01790_ _01799_ VPWR VGND _01804_ sg13g2_nor3_1
X_08050_ _01784_ _01785_ _01800_ _01803_ _01804_ VPWR 
+ VGND
+ _01805_ sg13g2_a221oi_1
X_08051_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ _01786_ _01805_ VPWR VGND _01806_ sg13g2_nor3_1
X_08052_ _01786_ _01805_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ VPWR VGND _01807_ sg13g2_o21ai_1
X_08053_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[5]\ VPWR VGND _01808_ sg13g2_buf_1
X_08054_ _01808_ VPWR VGND _01809_ sg13g2_buf_1
X_08055_ _01809_ VPWR VGND _01810_ sg13g2_buf_1
X_08056_ _01810_ _01782_ VPWR VGND _01811_ sg13g2_and2_1
X_08057_ _01739_ VPWR VGND _01812_ sg13g2_buf_1
X_08058_ _01734_ _01737_ VPWR VGND _01813_ sg13g2_xor2_1
X_08059_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[8]\ VPWR VGND _01814_ sg13g2_buf_1
X_08060_ _01758_ _01612_ _01616_ VPWR VGND _01815_ sg13g2_a21oi_1
X_08061_ _01753_ _01607_ VPWR VGND _01816_ sg13g2_xnor2_1
X_08062_ _01815_ _01816_ VPWR VGND _01817_ sg13g2_xnor2_1
X_08063_ _01764_ VPWR VGND _01818_ sg13g2_buf_1
X_08064_ _01818_ VPWR VGND _01819_ sg13g2_buf_1
X_08065_ _01759_ _01819_ _01762_ _01770_ VPWR VGND 
+ _01820_
+ sg13g2_nor4_1
X_08066_ _01770_ _01611_ VPWR VGND _01821_ sg13g2_nand2b_1
X_08067_ _01611_ _01770_ _01818_ VPWR VGND _01822_ sg13g2_nand3b_1
X_08068_ _01818_ _01821_ _01822_ VPWR VGND _01823_ sg13g2_o21ai_1
X_08069_ _01616_ _01823_ _01767_ VPWR VGND _01824_ sg13g2_mux2_1
X_08070_ _01820_ _01824_ _01757_ VPWR VGND _01825_ sg13g2_mux2_1
X_08071_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[6]\ VPWR VGND _01826_ sg13g2_buf_1
X_08072_ _01826_ VPWR VGND _01827_ sg13g2_buf_1
X_08073_ _01758_ _01762_ VPWR VGND _01828_ sg13g2_nand2_1
X_08074_ _01826_ _01765_ _01828_ VPWR VGND _01829_ sg13g2_nor3_1
X_08075_ _01815_ _01829_ VPWR VGND _01830_ sg13g2_or2_1
X_08076_ _01770_ _01826_ VPWR VGND _01831_ sg13g2_nand2b_1
X_08077_ _01764_ VPWR VGND _01832_ sg13g2_buf_1
X_08078_ _01762_ _01831_ _01832_ VPWR VGND _01833_ sg13g2_a21oi_1
X_08079_ _01826_ VPWR VGND _01834_ sg13g2_inv_1
X_08080_ _01834_ _01770_ _01762_ VPWR VGND _01835_ sg13g2_a21oi_1
X_08081_ _01833_ _01835_ _01780_ VPWR VGND _01836_ sg13g2_o21ai_1
X_08082_ _01818_ _01826_ VPWR VGND _01837_ sg13g2_nand2b_1
X_08083_ _01762_ _01770_ _01837_ VPWR VGND _01838_ sg13g2_nor3_1
X_08084_ _01757_ _01838_ VPWR VGND _01839_ sg13g2_nor2_1
X_08085_ _01760_ VPWR VGND _01840_ sg13g2_buf_1
X_08086_ _01840_ VPWR VGND _01841_ sg13g2_buf_1
X_08087_ _01757_ _01830_ _01836_ _01839_ _01841_ VPWR 
+ VGND
+ _01842_ sg13g2_a221oi_1
X_08088_ _01814_ _01817_ _01825_ _01827_ _01842_ VPWR 
+ VGND
+ _01843_ sg13g2_a221oi_1
X_08089_ _01812_ _01813_ _01843_ VPWR VGND _01844_ sg13g2_o21ai_1
X_08090_ _01782_ _01806_ _01807_ _01811_ _01844_ VPWR 
+ VGND
+ _01845_ sg13g2_a221oi_1
X_08091_ _01667_ _01633_ VPWR VGND _01846_ sg13g2_xor2_1
X_08092_ _01630_ _01631_ _01846_ VPWR VGND _01847_ sg13g2_nand3_1
X_08093_ _01630_ _01631_ _01846_ VPWR VGND _01848_ sg13g2_a21o_1
X_08094_ _00016_ VPWR VGND _01849_ sg13g2_buf_1
X_08095_ _01849_ VPWR VGND _01850_ sg13g2_buf_1
X_08096_ _01847_ _01848_ _01850_ VPWR VGND _01851_ sg13g2_a21o_1
X_08097_ _01752_ _01845_ _01851_ VPWR VGND _01852_ sg13g2_o21ai_1
X_08098_ _01717_ VPWR VGND _01853_ sg13g2_buf_1
X_08099_ _01849_ _01630_ _01631_ VPWR VGND _01854_ sg13g2_nand3_1
X_08100_ _01853_ _01633_ _01854_ VPWR VGND _01855_ sg13g2_nand3_1
X_08101_ _00015_ VPWR VGND _01856_ sg13g2_buf_1
X_08102_ _01661_ _01856_ VPWR VGND _01857_ sg13g2_xnor2_1
X_08103_ _01857_ VPWR VGND _01858_ sg13g2_buf_1
X_08104_ _01635_ _01858_ VPWR VGND _01859_ sg13g2_xor2_1
X_08105_ _01859_ _01847_ VPWR VGND _01860_ sg13g2_and2_1
X_08106_ _01717_ _01850_ _01665_ VPWR VGND _01861_ sg13g2_a21o_1
X_08107_ _01633_ _01630_ _01631_ VPWR VGND _01862_ sg13g2_nand3_1
X_08108_ _01717_ _01850_ VPWR VGND _01863_ sg13g2_nor2_1
X_08109_ _01862_ _01863_ _01859_ VPWR VGND _01864_ sg13g2_a21oi_1
X_08110_ _01855_ _01860_ _01861_ _01864_ VPWR VGND 
+ _01865_
+ sg13g2_a22oi_1
X_08111_ _01733_ _01852_ _01865_ VPWR VGND _01866_ sg13g2_o21ai_1
X_08112_ _01723_ _01726_ _01866_ VPWR VGND _01867_ sg13g2_o21ai_1
X_08113_ _01715_ _01716_ _01725_ VPWR VGND _01868_ sg13g2_a21o_1
X_08114_ _01710_ _01867_ _01868_ VPWR VGND _01869_ sg13g2_nand3b_1
X_08115_ _01703_ _01708_ _01869_ VPWR VGND _01870_ sg13g2_o21ai_1
X_08116_ _01672_ VPWR VGND _01871_ sg13g2_buf_1
X_08117_ _01871_ VPWR VGND _01872_ sg13g2_buf_1
X_08118_ _01872_ VPWR VGND _01873_ sg13g2_buf_1
X_08119_ _01598_ _01705_ _01873_ VPWR VGND _01874_ sg13g2_a21o_1
X_08120_ _01598_ _01705_ _01874_ VPWR VGND _01875_ sg13g2_o21ai_1
X_08121_ _01595_ VPWR VGND _01876_ sg13g2_buf_1
X_08122_ _01876_ VPWR VGND _01877_ sg13g2_buf_1
X_08123_ _01877_ _01596_ VPWR VGND _01878_ sg13g2_xnor2_1
X_08124_ _01875_ _01878_ VPWR VGND _01879_ sg13g2_xnor2_1
X_08125_ _00021_ VPWR VGND _01880_ sg13g2_buf_1
X_08126_ _01880_ VPWR VGND _01881_ sg13g2_buf_1
X_08127_ _01681_ _01593_ VPWR VGND _01882_ sg13g2_xor2_1
X_08128_ _01679_ _01882_ VPWR VGND _01883_ sg13g2_xnor2_1
X_08129_ _01881_ _01883_ VPWR VGND _01884_ sg13g2_xnor2_1
X_08130_ _01870_ _01879_ _01884_ VPWR VGND _01885_ sg13g2_o21ai_1
X_08131_ _00012_ VPWR VGND _01886_ sg13g2_inv_1
X_08132_ _01886_ VPWR VGND _01887_ sg13g2_buf_1
X_08133_ _01870_ _01879_ _01887_ VPWR VGND _01888_ sg13g2_a21oi_1
X_08134_ _01885_ _01888_ VPWR VGND _01889_ sg13g2_nor2_1
X_08135_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[16]\ VPWR VGND _01890_ sg13g2_buf_1
X_08136_ _01890_ _01883_ VPWR VGND _01891_ sg13g2_nand2_1
X_08137_ _01688_ _01891_ VPWR VGND _01892_ sg13g2_nand2_1
X_08138_ _01889_ _01892_ VPWR VGND _01893_ sg13g2_nor2_1
X_08139_ _01690_ VPWR VGND _01894_ sg13g2_inv_1
X_08140_ _01894_ VPWR VGND _01895_ sg13g2_buf_1
X_08141_ _01895_ _01891_ VPWR VGND _01896_ sg13g2_nand2_1
X_08142_ _01689_ VPWR VGND _01897_ sg13g2_buf_1
X_08143_ _01897_ _01688_ VPWR VGND _01898_ sg13g2_nand2_1
X_08144_ _01889_ _01896_ _01898_ VPWR VGND _01899_ sg13g2_o21ai_1
X_08145_ _01701_ _01893_ _01899_ VPWR VGND _01900_ sg13g2_nor3_1
X_08146_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2070_o[0]\ VPWR VGND _01901_ sg13g2_buf_1
X_08147_ _00949_ VPWR VGND _01902_ sg13g2_buf_1
X_08148_ _01902_ VPWR VGND _01903_ sg13g2_buf_1
X_08149_ _01901_ _01903_ VPWR VGND _01904_ sg13g2_nand2_1
X_08150_ _01900_ _01904_ _01244_ VPWR VGND _00431_ sg13g2_o21ai_1
X_08151_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[14]\ VPWR VGND _01905_ sg13g2_buf_1
X_08152_ _01671_ _01709_ VPWR VGND _01906_ sg13g2_xnor2_1
X_08153_ _01906_ VPWR VGND _01907_ sg13g2_buf_1
X_08154_ _01907_ VPWR VGND _01908_ sg13g2_buf_1
X_08155_ _01905_ _01908_ VPWR VGND _01909_ sg13g2_xor2_1
X_08156_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[13]\ VPWR VGND _01910_ sg13g2_buf_1
X_08157_ _01910_ VPWR VGND _01911_ sg13g2_inv_1
X_08158_ _01600_ VPWR VGND _01912_ sg13g2_buf_1
X_08159_ _01725_ VPWR VGND _01913_ sg13g2_buf_1
X_08160_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[12]\ VPWR VGND _01914_ sg13g2_buf_1
X_08161_ _01634_ VPWR VGND _01915_ sg13g2_inv_1
X_08162_ _01639_ VPWR VGND _01916_ sg13g2_inv_1
X_08163_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[9]\ VPWR VGND _01917_ sg13g2_buf_1
X_08164_ _01917_ VPWR VGND _01918_ sg13g2_inv_1
X_08165_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[7]\ VPWR VGND _01919_ sg13g2_buf_1
X_08166_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[6]\ VPWR VGND _01920_ sg13g2_buf_1
X_08167_ _01920_ _01764_ _01614_ VPWR VGND _01921_ sg13g2_a21o_1
X_08168_ _01758_ _01920_ _01764_ VPWR VGND _01922_ sg13g2_and3_1
X_08169_ _01919_ _01921_ _01922_ VPWR VGND _01923_ sg13g2_a21oi_1
X_08170_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[8]\ VPWR VGND _01924_ sg13g2_buf_1
X_08171_ _01924_ _01619_ VPWR VGND _01925_ sg13g2_nand2_1
X_08172_ _01924_ _01619_ VPWR VGND _01926_ sg13g2_nor2_1
X_08173_ _01918_ _01744_ _01923_ _01925_ _01926_ VPWR 
+ VGND
+ _01927_ sg13g2_a221oi_1
X_08174_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[10]\ VPWR VGND _01928_ sg13g2_buf_1
X_08175_ _01928_ _01627_ _01917_ _01603_ VPWR VGND 
+ _01929_
+ sg13g2_a22oi_1
X_08176_ _01929_ VPWR VGND _01930_ sg13g2_inv_1
X_08177_ _01928_ _01627_ VPWR VGND _01931_ sg13g2_or2_1
X_08178_ _01927_ _01930_ _01931_ VPWR VGND _01932_ sg13g2_o21ai_1
X_08179_ _01932_ VPWR VGND _01933_ sg13g2_buf_1
X_08180_ _01916_ _01933_ VPWR VGND _01934_ sg13g2_or2_1
X_08181_ _01934_ VPWR VGND _01935_ sg13g2_buf_1
X_08182_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[11]\ VPWR VGND _01936_ sg13g2_inv_1
X_08183_ _01916_ _01933_ _01936_ VPWR VGND _01937_ sg13g2_a21o_1
X_08184_ _01915_ _01935_ _01937_ VPWR VGND _01938_ sg13g2_nand3_1
X_08185_ _01935_ _01937_ _01915_ VPWR VGND _01939_ sg13g2_a21oi_1
X_08186_ _01914_ _01938_ _01939_ VPWR VGND _01940_ sg13g2_a21oi_1
X_08187_ _01911_ _01912_ _01913_ _01940_ VPWR VGND 
+ _01941_
+ sg13g2_nor4_1
X_08188_ _01910_ _01712_ VPWR VGND _01942_ sg13g2_nor2_1
X_08189_ _01910_ _01711_ _01914_ _01938_ _01939_ VPWR 
+ VGND
+ _01943_ sg13g2_a221oi_1
X_08190_ _01942_ _01943_ VPWR VGND _01944_ sg13g2_nor2_1
X_08191_ _01941_ _01944_ VPWR VGND _01945_ sg13g2_nand2b_1
X_08192_ _01713_ VPWR VGND _01946_ sg13g2_buf_1
X_08193_ _01946_ VPWR VGND _01947_ sg13g2_buf_1
X_08194_ _01910_ _01947_ VPWR VGND _01948_ sg13g2_xnor2_1
X_08195_ _01940_ _01948_ VPWR VGND _01949_ sg13g2_xnor2_1
X_08196_ _01935_ _01937_ VPWR VGND _01950_ sg13g2_nand2_1
X_08197_ _01719_ VPWR VGND _01951_ sg13g2_buf_1
X_08198_ _01914_ _01951_ VPWR VGND _01952_ sg13g2_xor2_1
X_08199_ _01950_ _01952_ VPWR VGND _01953_ sg13g2_xnor2_1
X_08200_ _01722_ VPWR VGND _01954_ sg13g2_buf_1
X_08201_ _01913_ _01949_ _01953_ _01954_ VPWR VGND 
+ _01955_
+ sg13g2_a22oi_1
X_08202_ _01841_ VPWR VGND _01956_ sg13g2_buf_1
X_08203_ _01832_ VPWR VGND _01957_ sg13g2_buf_1
X_08204_ _01920_ _01957_ VPWR VGND _01958_ sg13g2_nand2_1
X_08205_ _01759_ VPWR VGND _01959_ sg13g2_buf_1
X_08206_ _01919_ _01959_ VPWR VGND _01960_ sg13g2_xor2_1
X_08207_ _01958_ _01960_ VPWR VGND _01961_ sg13g2_xnor2_1
X_08208_ _01771_ VPWR VGND _01962_ sg13g2_inv_1
X_08209_ _01783_ VPWR VGND _01963_ sg13g2_inv_1
X_08210_ _01963_ VPWR VGND _01964_ sg13g2_buf_1
X_08211_ _01787_ VPWR VGND _01965_ sg13g2_inv_1
X_08212_ _01965_ VPWR VGND _01966_ sg13g2_buf_1
X_08213_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ _01966_ VPWR VGND _01967_ sg13g2_nand2_1
X_08214_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ _01788_ VPWR VGND _01968_ sg13g2_nand2b_1
X_08215_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ VPWR VGND _01969_ sg13g2_inv_1
X_08216_ _01791_ VPWR VGND _01970_ sg13g2_buf_1
X_08217_ _01969_ _01970_ _01795_ VPWR VGND _01971_ sg13g2_o21ai_1
X_08218_ _01795_ _01792_ VPWR VGND _01972_ sg13g2_nor2_1
X_08219_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ _01972_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ VPWR VGND _01973_ sg13g2_a21o_1
X_08220_ _01968_ _01971_ _01973_ VPWR VGND _01974_ sg13g2_nand3_1
X_08221_ _01803_ _01967_ _01974_ VPWR VGND _01975_ sg13g2_nand3_1
X_08222_ _01967_ _01974_ _01803_ VPWR VGND _01976_ sg13g2_a21oi_1
X_08223_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ _01964_ _01975_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ _01976_ VPWR 
+ VGND
+ _01977_ sg13g2_a221oi_1
X_08224_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _01809_ VPWR VGND _01978_ sg13g2_nand2b_1
X_08225_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ _01964_ _01978_ VPWR VGND _01979_ sg13g2_o21ai_1
X_08226_ _01808_ VPWR VGND _01980_ sg13g2_inv_1
X_08227_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _01980_ VPWR VGND _01981_ sg13g2_nand2_1
X_08228_ _01977_ _01979_ _01981_ VPWR VGND _01982_ sg13g2_o21ai_1
X_08229_ _01834_ VPWR VGND _01983_ sg13g2_buf_1
X_08230_ _01962_ _01982_ _01983_ VPWR VGND _01984_ sg13g2_o21ai_1
X_08231_ _01920_ _01957_ VPWR VGND _01985_ sg13g2_xor2_1
X_08232_ _01771_ _01982_ _01985_ VPWR VGND _01986_ sg13g2_o21ai_1
X_08233_ _01984_ _01985_ _01986_ VPWR VGND _01987_ sg13g2_o21ai_1
X_08234_ _01956_ _01961_ _01987_ VPWR VGND _01988_ sg13g2_o21ai_1
X_08235_ _01754_ VPWR VGND _01989_ sg13g2_inv_1
X_08236_ _01753_ VPWR VGND _01990_ sg13g2_buf_1
X_08237_ _01924_ _01990_ VPWR VGND _01991_ sg13g2_xnor2_1
X_08238_ _01923_ _01991_ VPWR VGND _01992_ sg13g2_xnor2_1
X_08239_ _01989_ _01992_ VPWR VGND _01993_ sg13g2_xnor2_1
X_08240_ _01956_ _01961_ _01993_ VPWR VGND _01994_ sg13g2_a21oi_1
X_08241_ _01923_ _01925_ _01926_ VPWR VGND _01995_ sg13g2_a21oi_1
X_08242_ _01917_ _01740_ VPWR VGND _01996_ sg13g2_xnor2_1
X_08243_ _01995_ _01996_ VPWR VGND _01997_ sg13g2_xnor2_1
X_08244_ _01814_ VPWR VGND _01998_ sg13g2_buf_1
X_08245_ _01998_ _01992_ VPWR VGND _01999_ sg13g2_nand2_1
X_08246_ _01997_ _01999_ VPWR VGND _02000_ sg13g2_nand2_1
X_08247_ _01812_ VPWR VGND _02001_ sg13g2_buf_1
X_08248_ _02001_ _01999_ VPWR VGND _02002_ sg13g2_nand2_1
X_08249_ _01988_ _01994_ _02000_ _02002_ VPWR VGND 
+ _02003_
+ sg13g2_a22oi_1
X_08250_ _01917_ _01740_ _01995_ VPWR VGND _02004_ sg13g2_a21o_1
X_08251_ _01917_ _01740_ _02004_ VPWR VGND _02005_ sg13g2_o21ai_1
X_08252_ _01928_ _02005_ VPWR VGND _02006_ sg13g2_xor2_1
X_08253_ _01750_ _02006_ VPWR VGND _02007_ sg13g2_xnor2_1
X_08254_ _02001_ _01997_ _02007_ VPWR VGND _02008_ sg13g2_a21oi_1
X_08255_ _02003_ _02008_ VPWR VGND _02009_ sg13g2_nor2b_1
X_08256_ _01730_ _02006_ VPWR VGND _02010_ sg13g2_xnor2_1
X_08257_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[11]\ _01853_ VPWR VGND _02011_ sg13g2_xnor2_1
X_08258_ _01933_ _02011_ VPWR VGND _02012_ sg13g2_nor2_1
X_08259_ _01933_ _02011_ VPWR VGND _02013_ sg13g2_and2_1
X_08260_ _01850_ VPWR VGND _02014_ sg13g2_inv_1
X_08261_ _02014_ VPWR VGND _02015_ sg13g2_buf_1
X_08262_ _02012_ _02013_ _02015_ VPWR VGND _02016_ sg13g2_o21ai_1
X_08263_ _01728_ _02010_ _02016_ VPWR VGND _02017_ sg13g2_o21ai_1
X_08264_ _01916_ VPWR VGND _02018_ sg13g2_buf_1
X_08265_ _02015_ _01933_ VPWR VGND _02019_ sg13g2_and2_1
X_08266_ _02014_ _01933_ VPWR VGND _02020_ sg13g2_nor2_1
X_08267_ _02014_ _01933_ VPWR VGND _02021_ sg13g2_nand2_1
X_08268_ _01853_ _02020_ _02021_ VPWR VGND _02022_ sg13g2_o21ai_1
X_08269_ _02018_ _02019_ _02022_ _01936_ VPWR VGND 
+ _02023_
+ sg13g2_a22oi_1
X_08270_ _01914_ _01858_ VPWR VGND _02024_ sg13g2_xnor2_1
X_08271_ _01936_ _02018_ _02020_ VPWR VGND _02025_ sg13g2_nor3_1
X_08272_ _02024_ _02012_ _02025_ VPWR VGND _02026_ sg13g2_nor3_1
X_08273_ _02023_ _02024_ _02026_ VPWR VGND _02027_ sg13g2_a21oi_1
X_08274_ _02009_ _02017_ _02027_ VPWR VGND _02028_ sg13g2_o21ai_1
X_08275_ _01724_ VPWR VGND _02029_ sg13g2_buf_1
X_08276_ _01946_ _02029_ VPWR VGND _02030_ sg13g2_nor2_1
X_08277_ _01912_ _01725_ VPWR VGND _02031_ sg13g2_nor2_1
X_08278_ _01600_ _01725_ VPWR VGND _02032_ sg13g2_nand2_1
X_08279_ _01910_ _02031_ _02032_ VPWR VGND _02033_ sg13g2_o21ai_1
X_08280_ _01911_ _02030_ _02033_ _01940_ _01909_ VPWR 
+ VGND
+ _02034_ sg13g2_a221oi_1
X_08281_ _01909_ _01945_ _01955_ _02028_ _02034_ VPWR 
+ VGND
+ _02035_ sg13g2_a221oi_1
X_08282_ _00012_ VPWR VGND _02036_ sg13g2_buf_1
X_08283_ _02036_ VPWR VGND _02037_ sg13g2_buf_1
X_08284_ _01905_ _01706_ VPWR VGND _02038_ sg13g2_or2_1
X_08285_ _01905_ _01672_ VPWR VGND _02039_ sg13g2_nand2_1
X_08286_ _01942_ _01943_ _02039_ VPWR VGND _02040_ sg13g2_o21ai_1
X_08287_ _02038_ _02040_ VPWR VGND _02041_ sg13g2_and2_1
X_08288_ _02041_ VPWR VGND _02042_ sg13g2_buf_1
X_08289_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[15]\ VPWR VGND _02043_ sg13g2_buf_1
X_08290_ _01877_ VPWR VGND _02044_ sg13g2_buf_1
X_08291_ _02043_ _02044_ VPWR VGND _02045_ sg13g2_xnor2_1
X_08292_ _02042_ _02045_ VPWR VGND _02046_ sg13g2_xnor2_1
X_08293_ _01702_ VPWR VGND _02047_ sg13g2_buf_1
X_08294_ _02047_ VPWR VGND _02048_ sg13g2_buf_1
X_08295_ _02048_ VPWR VGND _02049_ sg13g2_buf_1
X_08296_ _01872_ VPWR VGND _02050_ sg13g2_buf_1
X_08297_ _01905_ _02050_ VPWR VGND _02051_ sg13g2_xor2_1
X_08298_ _01944_ _02051_ VPWR VGND _02052_ sg13g2_xnor2_1
X_08299_ _02049_ _02052_ VPWR VGND _02053_ sg13g2_nand2_1
X_08300_ _02037_ _02046_ _02053_ VPWR VGND _02054_ sg13g2_o21ai_1
X_08301_ _02038_ _02040_ VPWR VGND _02055_ sg13g2_nand2_1
X_08302_ _02036_ _02042_ VPWR VGND _02056_ sg13g2_nand2_1
X_08303_ _02043_ _02044_ _02056_ VPWR VGND _02057_ sg13g2_nand3_1
X_08304_ _02055_ _02045_ _02057_ VPWR VGND _02058_ sg13g2_o21ai_1
X_08305_ _02036_ _02042_ VPWR VGND _02059_ sg13g2_nor2_1
X_08306_ _01674_ _02056_ _02059_ VPWR VGND _02060_ sg13g2_a21oi_1
X_08307_ _01674_ _01887_ _02055_ VPWR VGND _02061_ sg13g2_nand3_1
X_08308_ _02043_ _02060_ _02061_ VPWR VGND _02062_ sg13g2_o21ai_1
X_08309_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[16]\ VPWR VGND _02063_ sg13g2_buf_1
X_08310_ _01681_ VPWR VGND _02064_ sg13g2_buf_1
X_08311_ _02064_ _01880_ VPWR VGND _02065_ sg13g2_xnor2_1
X_08312_ _02063_ _02065_ VPWR VGND _02066_ sg13g2_xnor2_1
X_08313_ _02058_ _02062_ _02066_ VPWR VGND _02067_ sg13g2_mux2_1
X_08314_ _02035_ _02054_ _02067_ VPWR VGND _02068_ sg13g2_o21ai_1
X_08315_ _01890_ VPWR VGND _02069_ sg13g2_buf_1
X_08316_ _02043_ VPWR VGND _02070_ sg13g2_inv_1
X_08317_ _01674_ _02055_ _02070_ VPWR VGND _02071_ sg13g2_a21oi_1
X_08318_ _01877_ _02042_ _02071_ VPWR VGND _02072_ sg13g2_a21oi_1
X_08319_ _01682_ VPWR VGND _02073_ sg13g2_buf_1
X_08320_ _02063_ _02073_ VPWR VGND _02074_ sg13g2_xnor2_1
X_08321_ _02072_ _02074_ VPWR VGND _02075_ sg13g2_xnor2_1
X_08322_ _02069_ _02075_ VPWR VGND _02076_ sg13g2_nand2_1
X_08323_ _01689_ VPWR VGND _02077_ sg13g2_inv_1
X_08324_ _02063_ _01682_ VPWR VGND _02078_ sg13g2_nor2_1
X_08325_ _02063_ _01682_ VPWR VGND _02079_ sg13g2_nand2_1
X_08326_ _02072_ _02078_ _02079_ VPWR VGND _02080_ sg13g2_o21ai_1
X_08327_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[17]\ VPWR VGND _02081_ sg13g2_buf_1
X_08328_ _02081_ _01685_ VPWR VGND _02082_ sg13g2_xor2_1
X_08329_ _02080_ _02082_ VPWR VGND _02083_ sg13g2_xnor2_1
X_08330_ _02077_ _02083_ VPWR VGND _02084_ sg13g2_xnor2_1
X_08331_ _02068_ _02076_ _02084_ VPWR VGND _02085_ sg13g2_a21oi_1
X_08332_ _01690_ VPWR VGND _02086_ sg13g2_buf_1
X_08333_ _02086_ _02083_ VPWR VGND _02087_ sg13g2_and2_1
X_08334_ _01685_ VPWR VGND _02088_ sg13g2_buf_1
X_08335_ _02088_ VPWR VGND _02089_ sg13g2_buf_1
X_08336_ _02081_ _02089_ _02080_ VPWR VGND _02090_ sg13g2_o21ai_1
X_08337_ _02081_ _02089_ VPWR VGND _02091_ sg13g2_nand2_1
X_08338_ _02090_ _02091_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2087_o\ VPWR VGND _02092_ sg13g2_a21o_1
X_08339_ _02085_ _02087_ _02092_ VPWR VGND _02093_ sg13g2_o21ai_1
X_08340_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2085_o[0]\ VPWR VGND _02094_ sg13g2_buf_1
X_08341_ _02094_ VPWR VGND _02095_ sg13g2_inv_1
X_08342_ _01106_ VPWR VGND _02096_ sg13g2_buf_1
X_08343_ _02095_ _02096_ VPWR VGND _02097_ sg13g2_nor2_1
X_08344_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2082_o[0]\ VPWR VGND _02098_ sg13g2_buf_1
X_08345_ _02098_ VPWR VGND _02099_ sg13g2_inv_1
X_08346_ _02099_ _01903_ VPWR VGND _02100_ sg13g2_nor2_1
X_08347_ _02093_ _02097_ _02100_ VPWR VGND _00432_ sg13g2_a21o_1
X_08348_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2085_o[1]\ VPWR VGND _02101_ sg13g2_buf_1
X_08349_ _02101_ VPWR VGND _02102_ sg13g2_inv_1
X_08350_ _01106_ VPWR VGND _02103_ sg13g2_buf_1
X_08351_ _02102_ _02103_ VPWR VGND _02104_ sg13g2_nor2_1
X_08352_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2082_o[1]\ VPWR VGND _02105_ sg13g2_buf_1
X_08353_ _02105_ VPWR VGND _02106_ sg13g2_inv_1
X_08354_ _02106_ _01903_ VPWR VGND _02107_ sg13g2_nor2_1
X_08355_ _02093_ _02104_ _02107_ VPWR VGND _00433_ sg13g2_a21o_1
X_08356_ _01902_ VPWR VGND _02108_ sg13g2_buf_1
X_08357_ _02108_ VPWR VGND _02109_ sg13g2_buf_1
X_08358_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2088_o[0]\ VPWR VGND _02110_ sg13g2_buf_1
X_08359_ _02110_ VPWR VGND _02111_ sg13g2_buf_2
X_08360_ _02111_ VPWR VGND _02112_ sg13g2_inv_1
X_08361_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[17]\ VPWR VGND _02113_ sg13g2_buf_1
X_08362_ _02113_ VPWR VGND _02114_ sg13g2_inv_1
X_08363_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[14]\ VPWR VGND _02115_ sg13g2_buf_1
X_08364_ _01706_ _02115_ VPWR VGND _02116_ sg13g2_nand2_1
X_08365_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[13]\ VPWR VGND _02117_ sg13g2_buf_1
X_08366_ _02117_ VPWR VGND _02118_ sg13g2_inv_1
X_08367_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[12]\ VPWR VGND _02119_ sg13g2_buf_1
X_08368_ _02119_ VPWR VGND _02120_ sg13g2_inv_1
X_08369_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[11]\ VPWR VGND _02121_ sg13g2_inv_1
X_08370_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[10]\ VPWR VGND _02122_ sg13g2_buf_1
X_08371_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[8]\ VPWR VGND _02123_ sg13g2_buf_1
X_08372_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[6]\ VPWR VGND _02124_ sg13g2_buf_1
X_08373_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[7]\ VPWR VGND _02125_ sg13g2_buf_1
X_08374_ _01609_ _02124_ _02125_ VPWR VGND _02126_ sg13g2_a21o_1
X_08375_ _01609_ _02125_ _02124_ VPWR VGND _02127_ sg13g2_and3_1
X_08376_ _02127_ VPWR VGND _02128_ sg13g2_buf_1
X_08377_ _01605_ _02123_ _02126_ _01614_ _02128_ VPWR 
+ VGND
+ _02129_ sg13g2_a221oi_1
X_08378_ _01606_ _02123_ VPWR VGND _02130_ sg13g2_nor2_1
X_08379_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[9]\ VPWR VGND _02131_ sg13g2_inv_1
X_08380_ _02129_ _02130_ _02131_ VPWR VGND _02132_ sg13g2_o21ai_1
X_08381_ _02131_ _02129_ _02130_ VPWR VGND _02133_ sg13g2_nor3_1
X_08382_ _01604_ _02132_ _02133_ VPWR VGND _02134_ sg13g2_a21o_1
X_08383_ _02134_ VPWR VGND _02135_ sg13g2_buf_1
X_08384_ _02122_ _02135_ VPWR VGND _02136_ sg13g2_nand2_1
X_08385_ _02122_ _02135_ _01648_ VPWR VGND _02137_ sg13g2_o21ai_1
X_08386_ _02121_ _02136_ _02137_ VPWR VGND _02138_ sg13g2_nand3_1
X_08387_ _02136_ _02137_ _02121_ VPWR VGND _02139_ sg13g2_a21oi_1
X_08388_ _01666_ _02138_ _02139_ VPWR VGND _02140_ sg13g2_a21oi_1
X_08389_ _01600_ _02118_ _02120_ _01915_ _02140_ VPWR 
+ VGND
+ _02141_ sg13g2_a221oi_1
X_08390_ _02141_ VPWR VGND _02142_ sg13g2_buf_1
X_08391_ _01711_ _02117_ VPWR VGND _02143_ sg13g2_nand2_1
X_08392_ _01662_ _02117_ _02119_ VPWR VGND _02144_ sg13g2_nand3_1
X_08393_ _01711_ _01661_ _02119_ VPWR VGND _02145_ sg13g2_nand3_1
X_08394_ _02143_ _02144_ _02145_ VPWR VGND _02146_ sg13g2_nand3_1
X_08395_ _02146_ VPWR VGND _02147_ sg13g2_buf_1
X_08396_ _02142_ _02147_ VPWR VGND _02148_ sg13g2_nor2_1
X_08397_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[15]\ VPWR VGND _02149_ sg13g2_buf_1
X_08398_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[16]\ VPWR VGND _02150_ sg13g2_buf_1
X_08399_ _02149_ _02150_ VPWR VGND _02151_ sg13g2_nand2_1
X_08400_ _01595_ _02150_ VPWR VGND _02152_ sg13g2_nand2_1
X_08401_ _01706_ _02115_ VPWR VGND _02153_ sg13g2_nor2_1
X_08402_ _02153_ VPWR VGND _02154_ sg13g2_buf_1
X_08403_ _02116_ _02148_ _02151_ _02152_ _02154_ VPWR 
+ VGND
+ _02155_ sg13g2_a221oi_1
X_08404_ _01680_ _02149_ VPWR VGND _02156_ sg13g2_nand2_1
X_08405_ _01595_ _01680_ VPWR VGND _02157_ sg13g2_nand2_1
X_08406_ _02116_ _02148_ _02156_ _02157_ _02154_ VPWR 
+ VGND
+ _02158_ sg13g2_a221oi_1
X_08407_ _01680_ _02150_ VPWR VGND _02159_ sg13g2_nand2_1
X_08408_ _01595_ _02149_ _02150_ VPWR VGND _02160_ sg13g2_nand3_1
X_08409_ _01595_ _01680_ _02149_ VPWR VGND _02161_ sg13g2_nand3_1
X_08410_ _02159_ _02160_ _02161_ VPWR VGND _02162_ sg13g2_nand3_1
X_08411_ _02155_ _02158_ _02162_ VPWR VGND _02163_ sg13g2_or3_1
X_08412_ _02163_ VPWR VGND _02164_ sg13g2_buf_1
X_08413_ _02114_ _02164_ VPWR VGND _02165_ sg13g2_xnor2_1
X_08414_ _02113_ _02164_ VPWR VGND _02166_ sg13g2_and2_1
X_08415_ _02165_ _02166_ _01696_ VPWR VGND _02167_ sg13g2_mux2_1
X_08416_ _02113_ _02164_ VPWR VGND _02168_ sg13g2_nor2_1
X_08417_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2090_o\ _02167_ _02168_ _01697_ VPWR VGND 
+ _02169_
+ sg13g2_a22oi_1
X_08418_ _01895_ _02169_ VPWR VGND _02170_ sg13g2_nor2_1
X_08419_ _01667_ _02138_ _02139_ VPWR VGND _02171_ sg13g2_a21o_1
X_08420_ _02119_ _02171_ VPWR VGND _02172_ sg13g2_nand2_1
X_08421_ _02119_ _02171_ _01719_ VPWR VGND _02173_ sg13g2_o21ai_1
X_08422_ _02173_ VPWR VGND _02174_ sg13g2_buf_1
X_08423_ _01912_ _02029_ VPWR VGND _02175_ sg13g2_nor2_1
X_08424_ _02118_ _02175_ VPWR VGND _02176_ sg13g2_nand2_1
X_08425_ _02117_ _02030_ VPWR VGND _02177_ sg13g2_nand2_1
X_08426_ _02115_ _01907_ VPWR VGND _02178_ sg13g2_xnor2_1
X_08427_ _02172_ _02174_ _02176_ _02177_ _02178_ VPWR 
+ VGND
+ _02179_ sg13g2_a221oi_1
X_08428_ _02115_ _01908_ VPWR VGND _02180_ sg13g2_xor2_1
X_08429_ _02117_ _02180_ _02175_ VPWR VGND _02181_ sg13g2_nand3_1
X_08430_ _02118_ _02030_ _02178_ VPWR VGND _02182_ sg13g2_nand3_1
X_08431_ _02172_ _02174_ VPWR VGND _02183_ sg13g2_nand2_1
X_08432_ _02181_ _02182_ _02183_ VPWR VGND _02184_ sg13g2_a21oi_1
X_08433_ _01672_ _02115_ VPWR VGND _02185_ sg13g2_and2_1
X_08434_ _02185_ VPWR VGND _02186_ sg13g2_buf_1
X_08435_ _01703_ _02154_ _02186_ _02148_ VPWR VGND 
+ _02187_
+ sg13g2_nor4_1
X_08436_ _02154_ _02186_ _02047_ VPWR VGND _02188_ sg13g2_o21ai_1
X_08437_ _02142_ _02147_ _02188_ VPWR VGND _02189_ sg13g2_nor3_1
X_08438_ _02179_ _02184_ _02187_ _02189_ VPWR VGND 
+ _02190_
+ sg13g2_or4_1
X_08439_ _02186_ _02142_ _02147_ VPWR VGND _02191_ sg13g2_nor3_1
X_08440_ _02154_ _02191_ VPWR VGND _02192_ sg13g2_nor2_1
X_08441_ _01877_ _02149_ VPWR VGND _02193_ sg13g2_xnor2_1
X_08442_ _02192_ _02193_ VPWR VGND _02194_ sg13g2_xnor2_1
X_08443_ _02190_ _02194_ VPWR VGND _02195_ sg13g2_nor2b_1
X_08444_ _01887_ _02190_ VPWR VGND _02196_ sg13g2_nor2_1
X_08445_ _01748_ VPWR VGND _02197_ sg13g2_buf_1
X_08446_ _01764_ _02124_ VPWR VGND _02198_ sg13g2_nand2_1
X_08447_ _02125_ _02198_ VPWR VGND _02199_ sg13g2_xor2_1
X_08448_ _01759_ _02199_ VPWR VGND _02200_ sg13g2_xnor2_1
X_08449_ _01841_ _01989_ _02200_ VPWR VGND _02201_ sg13g2_nor3_1
X_08450_ _01759_ _02126_ _02128_ VPWR VGND _02202_ sg13g2_a21oi_1
X_08451_ _01753_ _02123_ VPWR VGND _02203_ sg13g2_xnor2_1
X_08452_ _02202_ _02203_ VPWR VGND _02204_ sg13g2_xnor2_1
X_08453_ _01814_ _02201_ _02204_ VPWR VGND _02205_ sg13g2_o21ai_1
X_08454_ _01956_ _01754_ _02200_ _02204_ VPWR VGND 
+ _02206_
+ sg13g2_or4_1
X_08455_ _01759_ _01840_ VPWR VGND _02207_ sg13g2_xnor2_1
X_08456_ _02123_ _01756_ VPWR VGND _02208_ sg13g2_xor2_1
X_08457_ _02126_ _02208_ VPWR VGND _02209_ sg13g2_nor2_1
X_08458_ _02128_ _02208_ _02209_ VPWR VGND _02210_ sg13g2_a21oi_1
X_08459_ _02207_ _02210_ VPWR VGND _02211_ sg13g2_nor2_1
X_08460_ _01959_ _01841_ _02208_ VPWR VGND _02212_ sg13g2_nand3_1
X_08461_ _01761_ VPWR VGND _02213_ sg13g2_inv_1
X_08462_ _02208_ _02213_ _01780_ VPWR VGND _02214_ sg13g2_nand3b_1
X_08463_ _02212_ _02214_ _02199_ VPWR VGND _02215_ sg13g2_a21oi_1
X_08464_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[115]\ VPWR VGND _02216_ sg13g2_inv_1
X_08465_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ VPWR VGND _02217_ sg13g2_nand2b_1
X_08466_ _02216_ _02217_ _01795_ VPWR VGND _02218_ sg13g2_o21ai_1
X_08467_ _02216_ _02217_ VPWR VGND _02219_ sg13g2_nand2_1
X_08468_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _02218_ _02219_ VPWR VGND 
+ _02220_
+ sg13g2_a22oi_1
X_08469_ _01801_ VPWR VGND _02221_ sg13g2_inv_1
X_08470_ _02221_ VPWR VGND _02222_ sg13g2_buf_1
X_08471_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ VPWR VGND _02223_ sg13g2_nor2_1
X_08472_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ VPWR VGND _02224_ sg13g2_nor2_1
X_08473_ _01963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ VPWR VGND _02225_ sg13g2_nor2_1
X_08474_ _02220_ _02223_ _02224_ _02225_ VPWR VGND 
+ _02226_
+ sg13g2_or4_1
X_08475_ _02124_ _01773_ VPWR VGND _02227_ sg13g2_xor2_1
X_08476_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ _01963_ VPWR VGND 
+ _02228_
+ sg13g2_a22oi_1
X_08477_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[119]\ VPWR VGND _02229_ sg13g2_buf_1
X_08478_ _01809_ _02229_ VPWR VGND _02230_ sg13g2_xnor2_1
X_08479_ _02225_ _02228_ _02230_ VPWR VGND _02231_ sg13g2_o21ai_1
X_08480_ _02227_ _02231_ VPWR VGND _02232_ sg13g2_nor2_1
X_08481_ _01771_ _01808_ VPWR VGND _02233_ sg13g2_nand2_1
X_08482_ _02233_ VPWR VGND _02234_ sg13g2_buf_1
X_08483_ _02229_ _02234_ _01983_ VPWR VGND _02235_ sg13g2_o21ai_1
X_08484_ _01818_ _02124_ VPWR VGND _02236_ sg13g2_xnor2_1
X_08485_ _01962_ _01809_ VPWR VGND _02237_ sg13g2_nand2_1
X_08486_ _02237_ VPWR VGND _02238_ sg13g2_buf_1
X_08487_ _02229_ _02236_ _02238_ VPWR VGND _02239_ sg13g2_nor3_1
X_08488_ _02235_ _02236_ _02239_ VPWR VGND _02240_ sg13g2_a21o_1
X_08489_ _02226_ _02232_ _02240_ VPWR VGND _02241_ sg13g2_a21o_1
X_08490_ _02211_ _02215_ _02241_ VPWR VGND _02242_ sg13g2_o21ai_1
X_08491_ _01812_ _02205_ _02206_ _02242_ VPWR VGND 
+ _02243_
+ sg13g2_nand4_1
X_08492_ _02129_ _02130_ VPWR VGND _02244_ sg13g2_nor2_1
X_08493_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[9]\ VPWR VGND _02245_ sg13g2_xnor2_1
X_08494_ _02244_ _02245_ VPWR VGND _02246_ sg13g2_xnor2_1
X_08495_ _02205_ _02206_ _02242_ _02246_ VPWR VGND 
+ _02247_
+ sg13g2_nand4_1
X_08496_ _01812_ _02246_ VPWR VGND _02248_ sg13g2_nand2_1
X_08497_ _02197_ _02243_ _02247_ _02248_ VPWR VGND 
+ _02249_
+ sg13g2_nand4_1
X_08498_ _01727_ VPWR VGND _02250_ sg13g2_buf_1
X_08499_ _01730_ _02122_ VPWR VGND _02251_ sg13g2_xnor2_1
X_08500_ _02135_ _02251_ VPWR VGND _02252_ sg13g2_xnor2_1
X_08501_ _02250_ _02252_ VPWR VGND _02253_ sg13g2_nor2_1
X_08502_ _01748_ VPWR VGND _02254_ sg13g2_inv_1
X_08503_ _02254_ _02243_ _02247_ _02248_ VPWR VGND 
+ _02255_
+ sg13g2_nand4_1
X_08504_ _02249_ _02253_ _02255_ _02252_ VPWR VGND 
+ _02256_
+ sg13g2_a22oi_1
X_08505_ _02136_ _02137_ VPWR VGND _02257_ sg13g2_nand2_1
X_08506_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[11]\ VPWR VGND _02258_ sg13g2_xor2_1
X_08507_ _02257_ _02258_ VPWR VGND _02259_ sg13g2_xnor2_1
X_08508_ _02015_ _02256_ _02259_ VPWR VGND _02260_ sg13g2_a21oi_1
X_08509_ _01719_ _02119_ VPWR VGND _02261_ sg13g2_xnor2_1
X_08510_ _02140_ _02261_ VPWR VGND _02262_ sg13g2_xnor2_1
X_08511_ _01856_ _02262_ VPWR VGND _02263_ sg13g2_xnor2_1
X_08512_ _02015_ _02256_ _02263_ VPWR VGND _02264_ sg13g2_o21ai_1
X_08513_ _01954_ _02262_ VPWR VGND _02265_ sg13g2_nand2_1
X_08514_ _02260_ _02264_ _02265_ VPWR VGND _02266_ sg13g2_o21ai_1
X_08515_ _02172_ _02174_ _02118_ VPWR VGND _02267_ sg13g2_a21oi_1
X_08516_ _02031_ _02267_ _02148_ VPWR VGND _02268_ sg13g2_a21oi_1
X_08517_ _02178_ _02268_ VPWR VGND _02269_ sg13g2_or2_1
X_08518_ _01725_ _02118_ _02172_ _02174_ VPWR VGND 
+ _02270_
+ sg13g2_nand4_1
X_08519_ _02032_ _02267_ _02270_ VPWR VGND _02271_ sg13g2_o21ai_1
X_08520_ _01947_ _02117_ _02183_ VPWR VGND _02272_ sg13g2_nor3_1
X_08521_ _02180_ _02271_ _02272_ VPWR VGND _02273_ sg13g2_or3_1
X_08522_ _02266_ _02269_ _02273_ VPWR VGND _02274_ sg13g2_nand3_1
X_08523_ _02195_ _02196_ _02274_ VPWR VGND _02275_ sg13g2_o21ai_1
X_08524_ _02037_ VPWR VGND _02276_ sg13g2_buf_1
X_08525_ _02276_ _02194_ VPWR VGND _02277_ sg13g2_nand2_1
X_08526_ _01881_ VPWR VGND _02278_ sg13g2_buf_1
X_08527_ _02149_ VPWR VGND _02279_ sg13g2_inv_1
X_08528_ _02279_ _02154_ _02191_ VPWR VGND _02280_ sg13g2_nor3_1
X_08529_ _02154_ _02191_ _02279_ VPWR VGND _02281_ sg13g2_o21ai_1
X_08530_ _02044_ _02280_ _02281_ VPWR VGND _02282_ sg13g2_o21ai_1
X_08531_ _01682_ _02150_ VPWR VGND _02283_ sg13g2_xnor2_1
X_08532_ _02282_ _02283_ VPWR VGND _02284_ sg13g2_xnor2_1
X_08533_ _02278_ _02284_ VPWR VGND _02285_ sg13g2_xnor2_1
X_08534_ _02275_ _02277_ _02285_ VPWR VGND _02286_ sg13g2_nand3_1
X_08535_ _02069_ _02284_ VPWR VGND _02287_ sg13g2_nand2_1
X_08536_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2090_o\ _01105_ VPWR VGND _02288_ sg13g2_nor2_1
X_08537_ _01686_ _01689_ VPWR VGND _02289_ sg13g2_nand2_1
X_08538_ _01696_ _02077_ VPWR VGND _02290_ sg13g2_nand2_1
X_08539_ _02288_ _02289_ _02290_ VPWR VGND _02291_ sg13g2_o21ai_1
X_08540_ _01686_ _01689_ VPWR VGND _02292_ sg13g2_xor2_1
X_08541_ _02288_ _02164_ _02113_ VPWR VGND _02293_ sg13g2_nand3b_1
X_08542_ _02113_ _02164_ _02293_ VPWR VGND _02294_ sg13g2_o21ai_1
X_08543_ _02165_ _02291_ _02292_ _02294_ VPWR VGND 
+ _02295_
+ sg13g2_a22oi_1
X_08544_ _02286_ _02287_ _02295_ VPWR VGND _02296_ sg13g2_a21oi_1
X_08545_ _02112_ _01107_ _02170_ _02296_ VPWR VGND 
+ _02297_
+ sg13g2_or4_1
X_08546_ _02095_ _02109_ _02297_ VPWR VGND _00434_ sg13g2_o21ai_1
X_08547_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2088_o[1]\ VPWR VGND _02298_ sg13g2_buf_1
X_08548_ _02298_ VPWR VGND _02299_ sg13g2_buf_2
X_08549_ _02299_ VPWR VGND _02300_ sg13g2_inv_1
X_08550_ _02300_ _01107_ _02170_ _02296_ VPWR VGND 
+ _02301_
+ sg13g2_or4_1
X_08551_ _02102_ _02109_ _02301_ VPWR VGND _00435_ sg13g2_o21ai_1
X_08552_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2091_o[0]\ VPWR VGND _02302_ sg13g2_buf_1
X_08553_ _02302_ VPWR VGND _02303_ sg13g2_inv_1
X_08554_ _01689_ _00949_ VPWR VGND _02304_ sg13g2_nand2_1
X_08555_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[12]\ VPWR VGND _02305_ sg13g2_inv_1
X_08556_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[11]\ VPWR VGND _02306_ sg13g2_inv_1
X_08557_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[10]\ VPWR VGND _02307_ sg13g2_buf_1
X_08558_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[8]\ VPWR VGND _02308_ sg13g2_buf_1
X_08559_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[6]\ VPWR VGND _02309_ sg13g2_buf_1
X_08560_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[7]\ VPWR VGND _02310_ sg13g2_buf_1
X_08561_ _01763_ _02309_ _02310_ VPWR VGND _02311_ sg13g2_a21o_1
X_08562_ _02311_ VPWR VGND _02312_ sg13g2_buf_1
X_08563_ _01764_ _02310_ _02309_ VPWR VGND _02313_ sg13g2_and3_1
X_08564_ _02313_ VPWR VGND _02314_ sg13g2_buf_1
X_08565_ _01619_ _02308_ _02312_ _01758_ _02314_ VPWR 
+ VGND
+ _02315_ sg13g2_a221oi_1
X_08566_ _01753_ _02308_ VPWR VGND _02316_ sg13g2_nor2_1
X_08567_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[9]\ VPWR VGND _02317_ sg13g2_inv_1
X_08568_ _02315_ _02316_ _02317_ VPWR VGND _02318_ sg13g2_o21ai_1
X_08569_ _02317_ _02315_ _02316_ VPWR VGND _02319_ sg13g2_nor3_1
X_08570_ _01735_ _02318_ _02319_ VPWR VGND _02320_ sg13g2_a21o_1
X_08571_ _02320_ VPWR VGND _02321_ sg13g2_buf_1
X_08572_ _02307_ _02321_ VPWR VGND _02322_ sg13g2_nand2_1
X_08573_ _02307_ _02321_ _01729_ VPWR VGND _02323_ sg13g2_o21ai_1
X_08574_ _02306_ _02322_ _02323_ VPWR VGND _02324_ sg13g2_nand3_1
X_08575_ _02322_ _02323_ _02306_ VPWR VGND _02325_ sg13g2_a21oi_1
X_08576_ _01717_ _02324_ _02325_ VPWR VGND _02326_ sg13g2_a21oi_1
X_08577_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[13]\ VPWR VGND _02327_ sg13g2_buf_1
X_08578_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[14]\ VPWR VGND _02328_ sg13g2_buf_1
X_08579_ _01713_ _02327_ _02328_ VPWR VGND _02329_ sg13g2_o21ai_1
X_08580_ _01713_ _02327_ _01706_ VPWR VGND _02330_ sg13g2_o21ai_1
X_08581_ _01667_ _02324_ _02325_ VPWR VGND _02331_ sg13g2_a21o_1
X_08582_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[12]\ _02331_ _01719_ VPWR VGND _02332_ sg13g2_a21oi_1
X_08583_ _02305_ _02326_ _02329_ _02330_ _02332_ VPWR 
+ VGND
+ _02333_ sg13g2_a221oi_1
X_08584_ _01675_ VPWR VGND _02334_ sg13g2_buf_1
X_08585_ _02328_ VPWR VGND _02335_ sg13g2_inv_1
X_08586_ _01713_ _02327_ VPWR VGND _02336_ sg13g2_nand2_1
X_08587_ _02334_ _02335_ _02336_ VPWR VGND _02337_ sg13g2_a21oi_1
X_08588_ _01871_ _02328_ _02337_ VPWR VGND _02338_ sg13g2_a21o_1
X_08589_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[15]\ VPWR VGND _02339_ sg13g2_buf_1
X_08590_ _02333_ _02338_ _02339_ VPWR VGND _02340_ sg13g2_o21ai_1
X_08591_ _02339_ _02333_ _02338_ VPWR VGND _02341_ sg13g2_nor3_1
X_08592_ _01674_ _02340_ _02341_ VPWR VGND _02342_ sg13g2_a21o_1
X_08593_ _02064_ VPWR VGND _02343_ sg13g2_buf_1
X_08594_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[16]\ VPWR VGND _02344_ sg13g2_buf_1
X_08595_ _02343_ _02344_ VPWR VGND _02345_ sg13g2_nand2_1
X_08596_ _02343_ _02344_ VPWR VGND _02346_ sg13g2_nor2_1
X_08597_ _02342_ _02345_ _02346_ VPWR VGND _02347_ sg13g2_a21oi_1
X_08598_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[17]\ VPWR VGND _02348_ sg13g2_buf_1
X_08599_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[17]\ _02348_ VPWR VGND _02349_ sg13g2_nor2_1
X_08600_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2093_o\ _02349_ _01690_ VPWR VGND _02350_ sg13g2_o21ai_1
X_08601_ _02350_ VPWR VGND _02351_ sg13g2_inv_1
X_08602_ _01689_ _01105_ _02351_ VPWR VGND _02352_ sg13g2_nor3_1
X_08603_ _02352_ _02347_ VPWR VGND _02353_ sg13g2_nor2_1
X_08604_ _02304_ _02347_ _02353_ VPWR VGND _02354_ sg13g2_a21oi_1
X_08605_ _02088_ _02348_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2093_o\ VPWR VGND _02355_ sg13g2_nand3_1
X_08606_ _02349_ _02355_ VPWR VGND _02356_ sg13g2_nand2b_1
X_08607_ _02354_ _02356_ VPWR VGND _02357_ sg13g2_nand2b_1
X_08608_ _02088_ _02348_ VPWR VGND _02358_ sg13g2_xor2_1
X_08609_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2093_o\ VPWR VGND _02359_ sg13g2_inv_1
X_08610_ _02359_ _02352_ VPWR VGND _02360_ sg13g2_nor2_1
X_08611_ _02304_ _02360_ _02347_ VPWR VGND _02361_ sg13g2_mux2_1
X_08612_ _02077_ _02351_ _02358_ _02361_ _01106_ VPWR 
+ VGND
+ _02362_ sg13g2_a221oi_1
X_08613_ _02305_ _02326_ _02332_ VPWR VGND _02363_ sg13g2_a21o_1
X_08614_ _01947_ _02327_ VPWR VGND _02364_ sg13g2_xnor2_1
X_08615_ _02363_ _02364_ VPWR VGND _02365_ sg13g2_xnor2_1
X_08616_ _02322_ _02323_ VPWR VGND _02366_ sg13g2_nand2_1
X_08617_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[11]\ VPWR VGND _02367_ sg13g2_xor2_1
X_08618_ _02366_ _02367_ VPWR VGND _02368_ sg13g2_xnor2_1
X_08619_ _02308_ _01756_ VPWR VGND _02369_ sg13g2_xor2_1
X_08620_ _01840_ _02314_ _02312_ VPWR VGND _02370_ sg13g2_o21ai_1
X_08621_ _01841_ _02312_ VPWR VGND _02371_ sg13g2_nor2_1
X_08622_ _01780_ _02370_ _02371_ VPWR VGND _02372_ sg13g2_a21oi_1
X_08623_ _01832_ _02309_ VPWR VGND _02373_ sg13g2_nand2_1
X_08624_ _01767_ _02310_ VPWR VGND _02374_ sg13g2_xnor2_1
X_08625_ _01832_ _01761_ _02309_ VPWR VGND _02375_ sg13g2_nand3_1
X_08626_ _01759_ _02310_ _02375_ VPWR VGND _02376_ sg13g2_nand3_1
X_08627_ _02373_ _02374_ _02376_ VPWR VGND _02377_ sg13g2_o21ai_1
X_08628_ _02377_ _02369_ VPWR VGND _02378_ sg13g2_nand2_1
X_08629_ _02369_ _02372_ _02378_ VPWR VGND _02379_ sg13g2_o21ai_1
X_08630_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ VPWR VGND _02380_ sg13g2_inv_1
X_08631_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ VPWR VGND _02381_ sg13g2_inv_1
X_08632_ _01788_ VPWR VGND _02382_ sg13g2_buf_1
X_08633_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ VPWR VGND _02383_ sg13g2_inv_1
X_08634_ _01970_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ VPWR VGND _02384_ sg13g2_nor2b_1
X_08635_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ _02384_ VPWR VGND _02385_ sg13g2_nand2_1
X_08636_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ _02384_ _01797_ VPWR VGND _02386_ sg13g2_o21ai_1
X_08637_ _02382_ _02383_ _02385_ _02386_ VPWR VGND 
+ _02387_
+ sg13g2_a22oi_1
X_08638_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ _01966_ _02387_ VPWR 
+ VGND
+ _02388_ sg13g2_a221oi_1
X_08639_ _01803_ _02380_ _02381_ _01784_ _02388_ VPWR 
+ VGND
+ _02389_ sg13g2_a221oi_1
X_08640_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[138]\ VPWR VGND _02390_ sg13g2_buf_1
X_08641_ _01980_ _02390_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ _01964_ VPWR VGND 
+ _02391_
+ sg13g2_a22oi_1
X_08642_ _02309_ _01774_ VPWR VGND _02392_ sg13g2_xnor2_1
X_08643_ _02391_ _02392_ VPWR VGND _02393_ sg13g2_nand2_1
X_08644_ _02390_ _02234_ _01983_ VPWR VGND _02394_ sg13g2_o21ai_1
X_08645_ _01832_ _02309_ VPWR VGND _02395_ sg13g2_xnor2_1
X_08646_ _02373_ _02374_ VPWR VGND _02396_ sg13g2_xnor2_1
X_08647_ _02390_ _02238_ _02395_ VPWR VGND _02397_ sg13g2_nor3_1
X_08648_ _02394_ _02395_ _02396_ _02213_ _02397_ VPWR 
+ VGND
+ _02398_ sg13g2_a221oi_1
X_08649_ _02389_ _02393_ _02398_ VPWR VGND _02399_ sg13g2_o21ai_1
X_08650_ _01959_ _02312_ _02314_ VPWR VGND _02400_ sg13g2_a21oi_1
X_08651_ _01990_ _02308_ VPWR VGND _02401_ sg13g2_xnor2_1
X_08652_ _02400_ _02401_ VPWR VGND _02402_ sg13g2_xnor2_1
X_08653_ _02379_ _02399_ _02402_ _01998_ VPWR VGND 
+ _02403_
+ sg13g2_a22oi_1
X_08654_ _02001_ _02403_ VPWR VGND _02404_ sg13g2_nor2_1
X_08655_ _02315_ _02316_ VPWR VGND _02405_ sg13g2_nor2_1
X_08656_ _01740_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[9]\ VPWR VGND _02406_ sg13g2_xnor2_1
X_08657_ _02405_ _02406_ VPWR VGND _02407_ sg13g2_xnor2_1
X_08658_ _02001_ _02403_ _02407_ VPWR VGND _02408_ sg13g2_a21oi_1
X_08659_ _02404_ _02408_ VPWR VGND _02409_ sg13g2_nor2_1
X_08660_ _01730_ _02307_ VPWR VGND _02410_ sg13g2_xnor2_1
X_08661_ _02321_ _02410_ VPWR VGND _02411_ sg13g2_xnor2_1
X_08662_ _02250_ _02411_ VPWR VGND _02412_ sg13g2_nor2_1
X_08663_ _02254_ _02409_ _02412_ VPWR VGND _02413_ sg13g2_o21ai_1
X_08664_ _02197_ _02409_ _02411_ VPWR VGND _02414_ sg13g2_o21ai_1
X_08665_ _02015_ _02368_ _02413_ _02414_ VPWR VGND 
+ _02415_
+ sg13g2_a22oi_1
X_08666_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[12]\ _02331_ VPWR VGND _02416_ sg13g2_xnor2_1
X_08667_ _01858_ _02416_ VPWR VGND _02417_ sg13g2_xor2_1
X_08668_ _02015_ _02368_ _02417_ VPWR VGND _02418_ sg13g2_o21ai_1
X_08669_ _01915_ VPWR VGND _02419_ sg13g2_buf_1
X_08670_ _02419_ _02416_ VPWR VGND _02420_ sg13g2_xnor2_1
X_08671_ _01954_ _02420_ VPWR VGND _02421_ sg13g2_nand2_1
X_08672_ _02415_ _02418_ _02421_ VPWR VGND _02422_ sg13g2_o21ai_1
X_08673_ _02365_ _02422_ _01913_ VPWR VGND _02423_ sg13g2_o21ai_1
X_08674_ _02365_ _02422_ VPWR VGND _02424_ sg13g2_nand2_1
X_08675_ _02333_ _02338_ VPWR VGND _02425_ sg13g2_nor2_1
X_08676_ _01877_ _02339_ VPWR VGND _02426_ sg13g2_xor2_1
X_08677_ _02425_ _02426_ VPWR VGND _02427_ sg13g2_xnor2_1
X_08678_ _01709_ VPWR VGND _02428_ sg13g2_buf_1
X_08679_ _01947_ _02327_ VPWR VGND _02429_ sg13g2_nor2_1
X_08680_ _02363_ _02336_ _02429_ VPWR VGND _02430_ sg13g2_a21oi_1
X_08681_ _01873_ _02328_ VPWR VGND _02431_ sg13g2_xor2_1
X_08682_ _02430_ _02431_ VPWR VGND _02432_ sg13g2_xnor2_1
X_08683_ _02428_ _02432_ VPWR VGND _02433_ sg13g2_xnor2_1
X_08684_ _02427_ _02433_ VPWR VGND _02434_ sg13g2_nand2b_1
X_08685_ _01887_ _02433_ VPWR VGND _02435_ sg13g2_nand2_1
X_08686_ _02423_ _02424_ _02434_ _02435_ VPWR VGND 
+ _02436_
+ sg13g2_a22oi_1
X_08687_ _02049_ _02432_ VPWR VGND _02437_ sg13g2_nand2_1
X_08688_ _02037_ _02427_ _02437_ VPWR VGND _02438_ sg13g2_a21o_1
X_08689_ _02276_ _02427_ _02438_ VPWR VGND _02439_ sg13g2_o21ai_1
X_08690_ _02073_ _02344_ VPWR VGND _02440_ sg13g2_xnor2_1
X_08691_ _02342_ _02440_ VPWR VGND _02441_ sg13g2_xnor2_1
X_08692_ _02278_ _02441_ VPWR VGND _02442_ sg13g2_xnor2_1
X_08693_ _02436_ _02439_ _02442_ VPWR VGND _02443_ sg13g2_o21ai_1
X_08694_ _02358_ _02347_ VPWR VGND _02444_ sg13g2_xnor2_1
X_08695_ _02069_ _02441_ _02444_ _02086_ _01106_ VPWR 
+ VGND
+ _02445_ sg13g2_a221oi_1
X_08696_ _02357_ _02362_ _02443_ _02445_ VPWR VGND 
+ _02446_
+ sg13g2_a22oi_1
X_08697_ _01106_ VPWR VGND _02447_ sg13g2_buf_1
X_08698_ _02447_ VPWR VGND _02448_ sg13g2_buf_1
X_08699_ _02111_ _02448_ VPWR VGND _02449_ sg13g2_nand2_1
X_08700_ _02303_ _02446_ _02449_ VPWR VGND _00436_ sg13g2_o21ai_1
X_08701_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2091_o[1]\ VPWR VGND _02450_ sg13g2_buf_1
X_08702_ _02450_ VPWR VGND _02451_ sg13g2_inv_1
X_08703_ _02299_ _02448_ VPWR VGND _02452_ sg13g2_nand2_1
X_08704_ _02451_ _02446_ _02452_ VPWR VGND _00437_ sg13g2_o21ai_1
X_08705_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[17]\ VPWR VGND _02453_ sg13g2_buf_1
X_08706_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[16]\ VPWR VGND _02454_ sg13g2_inv_1
X_08707_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[15]\ VPWR VGND _02455_ sg13g2_inv_1
X_08708_ _01674_ _02455_ VPWR VGND _02456_ sg13g2_nor2_1
X_08709_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[13]\ VPWR VGND _02457_ sg13g2_buf_1
X_08710_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[12]\ VPWR VGND _02458_ sg13g2_buf_1
X_08711_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[11]\ VPWR VGND _02459_ sg13g2_inv_1
X_08712_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[9]\ VPWR VGND _02460_ sg13g2_buf_1
X_08713_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[6]\ VPWR VGND _02461_ sg13g2_buf_1
X_08714_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[7]\ VPWR VGND _02462_ sg13g2_buf_1
X_08715_ _01609_ _02461_ _02462_ VPWR VGND _02463_ sg13g2_a21o_1
X_08716_ _01763_ _02462_ _02461_ VPWR VGND _02464_ sg13g2_and3_1
X_08717_ _01614_ _02463_ _02464_ VPWR VGND _02465_ sg13g2_a21oi_1
X_08718_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[8]\ VPWR VGND _02466_ sg13g2_buf_1
X_08719_ _01606_ _02466_ VPWR VGND _02467_ sg13g2_nand2_1
X_08720_ _01606_ _02466_ VPWR VGND _02468_ sg13g2_nor2_1
X_08721_ _02465_ _02467_ _02468_ VPWR VGND _02469_ sg13g2_a21oi_1
X_08722_ _01603_ _02460_ _02469_ VPWR VGND _02470_ sg13g2_o21ai_1
X_08723_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[10]\ VPWR VGND _02471_ sg13g2_buf_1
X_08724_ _01627_ _02471_ _02460_ _01603_ VPWR VGND 
+ _02472_
+ sg13g2_a22oi_1
X_08725_ _01627_ _02471_ VPWR VGND _02473_ sg13g2_nor2_1
X_08726_ _02470_ _02472_ _02473_ VPWR VGND _02474_ sg13g2_a21o_1
X_08727_ _02474_ VPWR VGND _02475_ sg13g2_buf_1
X_08728_ _02459_ _02475_ VPWR VGND _02476_ sg13g2_nor2_1
X_08729_ _02459_ _02475_ _01916_ VPWR VGND _02477_ sg13g2_a21oi_1
X_08730_ _02458_ _02476_ _02477_ VPWR VGND _02478_ sg13g2_nor3_1
X_08731_ _02476_ _02477_ _02458_ VPWR VGND _02479_ sg13g2_o21ai_1
X_08732_ _01915_ _02478_ _02479_ VPWR VGND _02480_ sg13g2_o21ai_1
X_08733_ _02457_ _02480_ VPWR VGND _02481_ sg13g2_nand2_1
X_08734_ _02457_ _02480_ _01713_ VPWR VGND _02482_ sg13g2_o21ai_1
X_08735_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[14]\ VPWR VGND _02483_ sg13g2_buf_1
X_08736_ _02483_ VPWR VGND _02484_ sg13g2_inv_1
X_08737_ _01674_ _02455_ _02481_ _02482_ _02484_ VPWR 
+ VGND
+ _02485_ sg13g2_a221oi_1
X_08738_ _01706_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[15]\ VPWR VGND _02486_ sg13g2_nand2_1
X_08739_ _01595_ _01706_ VPWR VGND _02487_ sg13g2_nand2_1
X_08740_ _02481_ _02482_ _02486_ _02487_ VPWR VGND 
+ _02488_
+ sg13g2_a22oi_1
X_08741_ _02486_ _02487_ _02484_ VPWR VGND _02489_ sg13g2_a21oi_1
X_08742_ _02456_ _02485_ _02488_ _02489_ VPWR VGND 
+ _02490_
+ sg13g2_nor4_1
X_08743_ _01681_ VPWR VGND _02491_ sg13g2_inv_1
X_08744_ _02454_ _02490_ _02491_ VPWR VGND _02492_ sg13g2_o21ai_1
X_08745_ _02454_ _02490_ VPWR VGND _02493_ sg13g2_nand2_1
X_08746_ _02492_ _02493_ VPWR VGND _02494_ sg13g2_and2_1
X_08747_ _02494_ VPWR VGND _02495_ sg13g2_buf_1
X_08748_ _02453_ _02495_ _02089_ VPWR VGND _02496_ sg13g2_o21ai_1
X_08749_ _02453_ _02495_ VPWR VGND _02497_ sg13g2_nand2_1
X_08750_ _02496_ _02497_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2096_o\ VPWR VGND _02498_ sg13g2_a21oi_1
X_08751_ _01686_ _02453_ VPWR VGND _02499_ sg13g2_xor2_1
X_08752_ _02495_ _02499_ VPWR VGND _02500_ sg13g2_xnor2_1
X_08753_ _01897_ _01691_ _02500_ VPWR VGND _02501_ sg13g2_mux2_1
X_08754_ _01107_ _02498_ _02501_ VPWR VGND _02502_ sg13g2_nor3_1
X_08755_ _02481_ _02482_ VPWR VGND _02503_ sg13g2_nand2_1
X_08756_ _02483_ _02503_ _02050_ VPWR VGND _02504_ sg13g2_a21o_1
X_08757_ _02483_ _02503_ _02504_ VPWR VGND _02505_ sg13g2_o21ai_1
X_08758_ _02044_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[15]\ VPWR VGND _02506_ sg13g2_xor2_1
X_08759_ _02505_ _02506_ VPWR VGND _02507_ sg13g2_xnor2_1
X_08760_ _02276_ _02507_ VPWR VGND _02508_ sg13g2_nand2_1
X_08761_ _01872_ _02483_ VPWR VGND _02509_ sg13g2_xor2_1
X_08762_ _02503_ _02509_ VPWR VGND _02510_ sg13g2_xnor2_1
X_08763_ _01946_ _02457_ VPWR VGND _02511_ sg13g2_xnor2_1
X_08764_ _02480_ _02511_ VPWR VGND _02512_ sg13g2_xnor2_1
X_08765_ _02512_ _01913_ VPWR VGND _02513_ sg13g2_nand2b_1
X_08766_ _02476_ _02477_ VPWR VGND _02514_ sg13g2_nor2_1
X_08767_ _01951_ _02458_ VPWR VGND _02515_ sg13g2_xnor2_1
X_08768_ _02514_ _02515_ VPWR VGND _02516_ sg13g2_xnor2_1
X_08769_ _01666_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[11]\ VPWR VGND _02517_ sg13g2_xor2_1
X_08770_ _02475_ _02517_ VPWR VGND _02518_ sg13g2_xnor2_1
X_08771_ _01849_ _02518_ VPWR VGND _02519_ sg13g2_nand2_1
X_08772_ _01735_ _02460_ VPWR VGND _02520_ sg13g2_xnor2_1
X_08773_ _02469_ _02520_ VPWR VGND _02521_ sg13g2_xnor2_1
X_08774_ _01738_ _02521_ VPWR VGND _02522_ sg13g2_nand2_1
X_08775_ _01753_ _02466_ VPWR VGND _02523_ sg13g2_xnor2_1
X_08776_ _02465_ _02523_ VPWR VGND _02524_ sg13g2_xnor2_1
X_08777_ _01754_ _02524_ VPWR VGND _02525_ sg13g2_nor2_1
X_08778_ _02522_ _02525_ VPWR VGND _02526_ sg13g2_and2_1
X_08779_ _01754_ _02522_ _02524_ VPWR VGND _02527_ sg13g2_and3_1
X_08780_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[157]\ VPWR VGND _02528_ sg13g2_buf_1
X_08781_ _02528_ _02234_ _01983_ VPWR VGND _02529_ sg13g2_o21ai_1
X_08782_ _01818_ _02461_ VPWR VGND _02530_ sg13g2_xnor2_1
X_08783_ _02528_ _02238_ _02530_ VPWR VGND _02531_ sg13g2_nor3_1
X_08784_ _02529_ _02530_ _02531_ VPWR VGND _02532_ sg13g2_a21o_1
X_08785_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ VPWR VGND _02533_ sg13g2_nor2b_1
X_08786_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _02533_ _01797_ VPWR VGND _02534_ sg13g2_a21oi_1
X_08787_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _02533_ VPWR VGND _02535_ sg13g2_nor2_1
X_08788_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[154]\ VPWR VGND _02536_ sg13g2_nand2_1
X_08789_ _02534_ _02535_ _02536_ VPWR VGND _02537_ sg13g2_o21ai_1
X_08790_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ VPWR VGND _02538_ sg13g2_inv_1
X_08791_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[154]\ VPWR VGND _02539_ sg13g2_inv_1
X_08792_ _01963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ VPWR VGND _02540_ sg13g2_nor2_1
X_08793_ _01802_ _02538_ _02539_ _01788_ _02540_ VPWR 
+ VGND
+ _02541_ sg13g2_a221oi_1
X_08794_ _02461_ _01773_ VPWR VGND _02542_ sg13g2_nand2_1
X_08795_ _02461_ _01773_ VPWR VGND _02543_ sg13g2_or2_1
X_08796_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ _01963_ VPWR VGND 
+ _02544_
+ sg13g2_a22oi_1
X_08797_ _01809_ _02528_ VPWR VGND _02545_ sg13g2_xnor2_1
X_08798_ _02540_ _02544_ _02545_ VPWR VGND _02546_ sg13g2_o21ai_1
X_08799_ _02537_ _02541_ _02542_ _02543_ _02546_ VPWR 
+ VGND
+ _02547_ sg13g2_a221oi_1
X_08800_ _02213_ VPWR VGND _02548_ sg13g2_buf_1
X_08801_ _02532_ _02547_ _02548_ VPWR VGND _02549_ sg13g2_o21ai_1
X_08802_ _01957_ _02461_ VPWR VGND _02550_ sg13g2_nand2_1
X_08803_ _01959_ _02462_ VPWR VGND _02551_ sg13g2_xor2_1
X_08804_ _02550_ _02551_ VPWR VGND _02552_ sg13g2_xnor2_1
X_08805_ _02548_ _02532_ _02547_ VPWR VGND _02553_ sg13g2_nor3_1
X_08806_ _02549_ _02552_ _02553_ VPWR VGND _02554_ sg13g2_a21oi_1
X_08807_ _02526_ _02527_ _02554_ VPWR VGND _02555_ sg13g2_o21ai_1
X_08808_ _01814_ _02524_ VPWR VGND _02556_ sg13g2_and2_1
X_08809_ _01812_ _02521_ VPWR VGND _02557_ sg13g2_nor2_1
X_08810_ _02522_ _02556_ _02557_ VPWR VGND _02558_ sg13g2_a21oi_1
X_08811_ _02460_ _02469_ _01736_ VPWR VGND _02559_ sg13g2_a21oi_1
X_08812_ _02460_ _02469_ VPWR VGND _02560_ sg13g2_nor2_1
X_08813_ _02559_ _02560_ VPWR VGND _02561_ sg13g2_nor2_1
X_08814_ _01729_ _02471_ VPWR VGND _02562_ sg13g2_xnor2_1
X_08815_ _02561_ _02562_ VPWR VGND _02563_ sg13g2_xnor2_1
X_08816_ _01748_ _02563_ VPWR VGND _02564_ sg13g2_xnor2_1
X_08817_ _02555_ _02558_ _02564_ VPWR VGND _02565_ sg13g2_a21oi_1
X_08818_ _01728_ _02563_ VPWR VGND _02566_ sg13g2_nor2_1
X_08819_ _01850_ _02518_ VPWR VGND _02567_ sg13g2_nor2_1
X_08820_ _02519_ _02566_ _02567_ VPWR VGND _02568_ sg13g2_a21o_1
X_08821_ _02519_ _02565_ _02568_ VPWR VGND _02569_ sg13g2_a21oi_1
X_08822_ _01856_ _02516_ _02569_ VPWR VGND _02570_ sg13g2_nor3_1
X_08823_ _01856_ VPWR VGND _02571_ sg13g2_inv_1
X_08824_ _01722_ VPWR VGND _02572_ sg13g2_inv_1
X_08825_ _02571_ _02569_ _02572_ VPWR VGND _02573_ sg13g2_o21ai_1
X_08826_ _02516_ _02573_ VPWR VGND _02574_ sg13g2_and2_1
X_08827_ _02029_ VPWR VGND _02575_ sg13g2_buf_1
X_08828_ _02575_ _02512_ VPWR VGND _02576_ sg13g2_nand2_1
X_08829_ _02570_ _02574_ _02576_ VPWR VGND _02577_ sg13g2_o21ai_1
X_08830_ _02428_ _02510_ VPWR VGND _02578_ sg13g2_or2_1
X_08831_ _02428_ _02510_ VPWR VGND _02579_ sg13g2_nand2_1
X_08832_ _02513_ _02577_ _02578_ _02579_ VPWR VGND 
+ _02580_
+ sg13g2_a22oi_1
X_08833_ _02049_ _02510_ _02580_ VPWR VGND _02581_ sg13g2_a21o_1
X_08834_ _02276_ _02507_ VPWR VGND _02582_ sg13g2_nor2_1
X_08835_ _02508_ _02581_ _02582_ VPWR VGND _02583_ sg13g2_a21oi_1
X_08836_ _02454_ _02490_ VPWR VGND _02584_ sg13g2_xnor2_1
X_08837_ _02065_ _02584_ VPWR VGND _02585_ sg13g2_xnor2_1
X_08838_ _02491_ _02584_ VPWR VGND _02586_ sg13g2_xnor2_1
X_08839_ _02086_ _02500_ _02586_ _02069_ VPWR VGND 
+ _02587_
+ sg13g2_a22oi_1
X_08840_ _02583_ _02585_ _02587_ VPWR VGND _02588_ sg13g2_o21ai_1
X_08841_ _01105_ VPWR VGND _02589_ sg13g2_buf_1
X_08842_ _02589_ VPWR VGND _02590_ sg13g2_buf_1
X_08843_ _02302_ _02590_ VPWR VGND _02591_ sg13g2_nand2_1
X_08844_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2094_o[0]\ VPWR VGND _02592_ sg13g2_buf_1
X_08845_ _01902_ VPWR VGND _02593_ sg13g2_buf_1
X_08846_ _02592_ _02593_ VPWR VGND _02594_ sg13g2_nand2_1
X_08847_ _02502_ _02588_ _02591_ _02594_ VPWR VGND 
+ _00438_
+ sg13g2_a22oi_1
X_08848_ _02450_ _02590_ VPWR VGND _02595_ sg13g2_nand2_1
X_08849_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2094_o[1]\ VPWR VGND _02596_ sg13g2_buf_1
X_08850_ _02596_ _02593_ VPWR VGND _02597_ sg13g2_nand2_1
X_08851_ _02502_ _02588_ _02595_ _02597_ VPWR VGND 
+ _00439_
+ sg13g2_a22oi_1
X_08852_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[15]\ VPWR VGND _02598_ sg13g2_buf_1
X_08853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[16]\ VPWR VGND _02599_ sg13g2_buf_1
X_08854_ _01877_ _02598_ _02599_ VPWR VGND _02600_ sg13g2_a21o_1
X_08855_ _01877_ _02598_ _01682_ VPWR VGND _02601_ sg13g2_a21o_1
X_08856_ _01876_ _02598_ VPWR VGND _02602_ sg13g2_nor2_1
X_08857_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[14]\ VPWR VGND _02603_ sg13g2_buf_1
X_08858_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[13]\ VPWR VGND _02604_ sg13g2_buf_1
X_08859_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[12]\ VPWR VGND _02605_ sg13g2_buf_1
X_08860_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[11]\ VPWR VGND _02606_ sg13g2_buf_1
X_08861_ _02606_ VPWR VGND _02607_ sg13g2_inv_1
X_08862_ _02018_ _02607_ VPWR VGND _02608_ sg13g2_nor2_1
X_08863_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[10]\ VPWR VGND _02609_ sg13g2_buf_1
X_08864_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[9]\ VPWR VGND _02610_ sg13g2_inv_1
X_08865_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[8]\ VPWR VGND _02611_ sg13g2_buf_1
X_08866_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[6]\ VPWR VGND _02612_ sg13g2_buf_1
X_08867_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[7]\ VPWR VGND _02613_ sg13g2_buf_1
X_08868_ _01609_ _02612_ _02613_ VPWR VGND _02614_ sg13g2_a21oi_1
X_08869_ _01763_ _02613_ _02612_ VPWR VGND _02615_ sg13g2_nand3_1
X_08870_ _01779_ _02614_ _02615_ VPWR VGND _02616_ sg13g2_o21ai_1
X_08871_ _02611_ _02616_ VPWR VGND _02617_ sg13g2_nand2_1
X_08872_ _02611_ _02616_ _01619_ VPWR VGND _02618_ sg13g2_o21ai_1
X_08873_ _02610_ _02617_ _02618_ VPWR VGND _02619_ sg13g2_nand3_1
X_08874_ _02617_ _02618_ _02610_ VPWR VGND _02620_ sg13g2_a21oi_1
X_08875_ _01604_ _02619_ _02620_ VPWR VGND _02621_ sg13g2_a21o_1
X_08876_ _02621_ VPWR VGND _02622_ sg13g2_buf_1
X_08877_ _02609_ _02622_ VPWR VGND _02623_ sg13g2_nand2_1
X_08878_ _02609_ _02622_ _01648_ VPWR VGND _02624_ sg13g2_o21ai_1
X_08879_ _02018_ _02607_ _02623_ _02624_ VPWR VGND 
+ _02625_
+ sg13g2_a22oi_1
X_08880_ _02625_ VPWR VGND _02626_ sg13g2_buf_1
X_08881_ _02604_ _02605_ _02608_ _02626_ VPWR VGND 
+ _02627_
+ sg13g2_nor4_1
X_08882_ _01711_ _02605_ _02608_ _02626_ VPWR VGND 
+ _02628_
+ sg13g2_nor4_1
X_08883_ _01661_ _02604_ VPWR VGND _02629_ sg13g2_or2_1
X_08884_ _01600_ _01915_ VPWR VGND _02630_ sg13g2_nand2_1
X_08885_ _01667_ _02606_ _02629_ _02630_ _02626_ VPWR 
+ VGND
+ _02631_ sg13g2_a221oi_1
X_08886_ _02629_ _02630_ _02605_ VPWR VGND _02632_ sg13g2_a21o_1
X_08887_ _01712_ _02604_ _02632_ VPWR VGND _02633_ sg13g2_o21ai_1
X_08888_ _02627_ _02628_ _02631_ _02633_ VPWR VGND 
+ _02634_
+ sg13g2_nor4_1
X_08889_ _02634_ VPWR VGND _02635_ sg13g2_buf_2
X_08890_ _02603_ _02635_ VPWR VGND _02636_ sg13g2_nor2_1
X_08891_ _02603_ _02635_ _01872_ VPWR VGND _02637_ sg13g2_a21oi_1
X_08892_ _02602_ _02636_ _02637_ VPWR VGND _02638_ sg13g2_nor3_1
X_08893_ _02600_ _02601_ _02638_ VPWR VGND _02639_ sg13g2_a21oi_1
X_08894_ _02343_ _02599_ VPWR VGND _02640_ sg13g2_nor2_1
X_08895_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[17]\ VPWR VGND _02641_ sg13g2_buf_1
X_08896_ _01685_ _02641_ VPWR VGND _02642_ sg13g2_xnor2_1
X_08897_ _02077_ _02639_ _02640_ _02642_ VPWR VGND 
+ _02643_
+ sg13g2_nor4_1
X_08898_ _02600_ _02601_ _02638_ VPWR VGND _02644_ sg13g2_a21o_1
X_08899_ _02073_ _02599_ VPWR VGND _02645_ sg13g2_or2_1
X_08900_ _02642_ VPWR VGND _02646_ sg13g2_inv_1
X_08901_ _02077_ _02646_ VPWR VGND _02647_ sg13g2_nand2_1
X_08902_ _02644_ _02645_ _02647_ VPWR VGND _02648_ sg13g2_a21oi_1
X_08903_ _01897_ _02639_ _02640_ _02646_ VPWR VGND 
+ _02649_
+ sg13g2_nor4_1
X_08904_ _01897_ _02642_ VPWR VGND _02650_ sg13g2_nand2_1
X_08905_ _02644_ _02645_ _02650_ VPWR VGND _02651_ sg13g2_a21oi_1
X_08906_ _02643_ _02648_ _02649_ _02651_ VPWR VGND 
+ _02652_
+ sg13g2_nor4_1
X_08907_ _01594_ _02598_ VPWR VGND _02653_ sg13g2_xor2_1
X_08908_ _02653_ VPWR VGND _02654_ sg13g2_buf_1
X_08909_ _02334_ _02636_ VPWR VGND _02655_ sg13g2_nand2_1
X_08910_ _02603_ _02635_ VPWR VGND _02656_ sg13g2_xnor2_1
X_08911_ _02050_ _02656_ _02637_ VPWR VGND _02657_ sg13g2_a21oi_1
X_08912_ _02654_ _02657_ VPWR VGND _02658_ sg13g2_nand2_1
X_08913_ _02654_ _02655_ _02658_ VPWR VGND _02659_ sg13g2_o21ai_1
X_08914_ _02605_ _02608_ _02626_ VPWR VGND _02660_ sg13g2_nor3_1
X_08915_ _02608_ _02626_ _02605_ VPWR VGND _02661_ sg13g2_o21ai_1
X_08916_ _02419_ _02660_ _02661_ VPWR VGND _02662_ sg13g2_o21ai_1
X_08917_ _01946_ _02604_ VPWR VGND _02663_ sg13g2_xnor2_1
X_08918_ _02662_ _02663_ VPWR VGND _02664_ sg13g2_xnor2_1
X_08919_ _02664_ _01913_ VPWR VGND _02665_ sg13g2_nand2b_1
X_08920_ _01871_ _02603_ VPWR VGND _02666_ sg13g2_xor2_1
X_08921_ _02635_ _02654_ _02666_ VPWR VGND _02667_ sg13g2_nand3b_1
X_08922_ _02603_ VPWR VGND _02668_ sg13g2_inv_1
X_08923_ _02334_ _02668_ _02635_ _02654_ VPWR VGND 
+ _02669_
+ sg13g2_nand4_1
X_08924_ _02047_ _02668_ _02654_ VPWR VGND _02670_ sg13g2_nor3_1
X_08925_ _02334_ _02668_ _02654_ VPWR VGND _02671_ sg13g2_nor3_1
X_08926_ _02670_ _02671_ _02635_ VPWR VGND _02672_ sg13g2_o21ai_1
X_08927_ _02334_ _02047_ _02653_ VPWR VGND _02673_ sg13g2_nor3_1
X_08928_ _01871_ _02047_ _02603_ VPWR VGND _02674_ sg13g2_nor3_1
X_08929_ _02334_ _02047_ _02668_ _02653_ VPWR VGND 
+ _02675_
+ sg13g2_nor4_1
X_08930_ _02635_ _02673_ _02674_ _02654_ _02675_ VPWR 
+ VGND
+ _02676_ sg13g2_a221oi_1
X_08931_ _02667_ _02669_ _02672_ _02676_ VPWR VGND 
+ _02677_
+ sg13g2_nand4_1
X_08932_ _01908_ _02656_ VPWR VGND _02678_ sg13g2_xnor2_1
X_08933_ _02677_ _02678_ _02037_ VPWR VGND _02679_ sg13g2_a21o_1
X_08934_ _02608_ _02626_ VPWR VGND _02680_ sg13g2_nor2_1
X_08935_ _01719_ _02605_ VPWR VGND _02681_ sg13g2_xnor2_1
X_08936_ _02680_ _02681_ VPWR VGND _02682_ sg13g2_xnor2_1
X_08937_ _01954_ _02682_ VPWR VGND _02683_ sg13g2_nand2_1
X_08938_ _02609_ _02622_ VPWR VGND _02684_ sg13g2_xnor2_1
X_08939_ _01628_ _02684_ VPWR VGND _02685_ sg13g2_xnor2_1
X_08940_ _01750_ _02684_ VPWR VGND _02686_ sg13g2_xor2_1
X_08941_ _01738_ VPWR VGND _02687_ sg13g2_inv_1
X_08942_ _02617_ _02618_ VPWR VGND _02688_ sg13g2_nand2_1
X_08943_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[9]\ VPWR VGND _02689_ sg13g2_xor2_1
X_08944_ _02688_ _02689_ VPWR VGND _02690_ sg13g2_xnor2_1
X_08945_ _02687_ _02690_ VPWR VGND _02691_ sg13g2_and2_1
X_08946_ _01727_ _02685_ _02686_ _02691_ VPWR VGND 
+ _02692_
+ sg13g2_a22oi_1
X_08947_ _01832_ _02612_ VPWR VGND _02693_ sg13g2_nand2_1
X_08948_ _01767_ _02613_ VPWR VGND _02694_ sg13g2_xnor2_1
X_08949_ _02693_ _02694_ VPWR VGND _02695_ sg13g2_xnor2_1
X_08950_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[176]\ VPWR VGND _02696_ sg13g2_buf_1
X_08951_ _02696_ _02234_ _01834_ VPWR VGND _02697_ sg13g2_o21ai_1
X_08952_ _01764_ _02612_ VPWR VGND _02698_ sg13g2_xor2_1
X_08953_ _02696_ _02238_ _02698_ VPWR VGND _02699_ sg13g2_o21ai_1
X_08954_ _02697_ _02698_ _02699_ VPWR VGND _02700_ sg13g2_o21ai_1
X_08955_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[172]\ VPWR VGND _02701_ sg13g2_inv_1
X_08956_ _01791_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ VPWR VGND _02702_ sg13g2_nand2b_1
X_08957_ _02701_ _02702_ VPWR VGND _02703_ sg13g2_nand2_1
X_08958_ _02701_ _02702_ VPWR VGND _02704_ sg13g2_nor2_1
X_08959_ _01965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _02703_ _01796_ _02704_ VPWR 
+ VGND
+ _02705_ sg13g2_a221oi_1
X_08960_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _01801_ VPWR VGND _02706_ sg13g2_nand2b_1
X_08961_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _01787_ VPWR VGND _02707_ sg13g2_nand2b_1
X_08962_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[4]\ VPWR VGND _02708_ sg13g2_nand2b_1
X_08963_ _02706_ _02707_ _02708_ VPWR VGND _02709_ sg13g2_nand3_1
X_08964_ _02612_ _01773_ VPWR VGND _02710_ sg13g2_xnor2_1
X_08965_ _01980_ _02696_ VPWR VGND _02711_ sg13g2_nand2_1
X_08966_ _02696_ VPWR VGND _02712_ sg13g2_inv_1
X_08967_ _01809_ _02712_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ _01963_ VPWR VGND 
+ _02713_
+ sg13g2_a22oi_1
X_08968_ _02221_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _02708_ VPWR VGND _02714_ sg13g2_nand3_1
X_08969_ _02710_ _02711_ _02713_ _02714_ VPWR VGND 
+ _02715_
+ sg13g2_and4_1
X_08970_ _02705_ _02709_ _02715_ VPWR VGND _02716_ sg13g2_o21ai_1
X_08971_ _01840_ _02700_ _02716_ VPWR VGND _02717_ sg13g2_nand3_1
X_08972_ _02700_ _02716_ _01841_ VPWR VGND _02718_ sg13g2_a21oi_1
X_08973_ _02695_ _02717_ _02718_ VPWR VGND _02719_ sg13g2_a21oi_1
X_08974_ _01753_ _02611_ VPWR VGND _02720_ sg13g2_xnor2_1
X_08975_ _02616_ _02720_ VPWR VGND _02721_ sg13g2_xnor2_1
X_08976_ _01814_ _02721_ VPWR VGND _02722_ sg13g2_nor2_1
X_08977_ _01989_ _02719_ _02722_ VPWR VGND _02723_ sg13g2_o21ai_1
X_08978_ _01754_ _02719_ _02721_ VPWR VGND _02724_ sg13g2_o21ai_1
X_08979_ _02686_ _02690_ _02723_ _02724_ VPWR VGND 
+ _02725_
+ sg13g2_nand4_1
X_08980_ _02687_ _02686_ _02723_ _02724_ VPWR VGND 
+ _02726_
+ sg13g2_nand4_1
X_08981_ _02692_ _02725_ _02726_ VPWR VGND _02727_ sg13g2_and3_1
X_08982_ _02623_ _02624_ VPWR VGND _02728_ sg13g2_nand2_1
X_08983_ _01717_ _02606_ VPWR VGND _02729_ sg13g2_xnor2_1
X_08984_ _02728_ _02729_ VPWR VGND _02730_ sg13g2_xnor2_1
X_08985_ _01849_ VPWR VGND _02731_ sg13g2_buf_1
X_08986_ _02727_ _02730_ _02731_ VPWR VGND _02732_ sg13g2_a21oi_1
X_08987_ _02727_ _02730_ VPWR VGND _02733_ sg13g2_nor2_1
X_08988_ _01856_ _02682_ VPWR VGND _02734_ sg13g2_xnor2_1
X_08989_ _02732_ _02733_ _02734_ VPWR VGND _02735_ sg13g2_o21ai_1
X_08990_ _02029_ _02664_ VPWR VGND _02736_ sg13g2_and2_1
X_08991_ _02683_ _02735_ _02736_ VPWR VGND _02737_ sg13g2_a21o_1
X_08992_ _02665_ _02679_ _02737_ VPWR VGND _02738_ sg13g2_nand3_1
X_08993_ _01908_ VPWR VGND _02739_ sg13g2_inv_1
X_08994_ _02603_ _02635_ VPWR VGND _02740_ sg13g2_and2_1
X_08995_ _02636_ _02740_ _02654_ VPWR VGND _02741_ sg13g2_mux2_1
X_08996_ _02050_ _02428_ _02654_ VPWR VGND _02742_ sg13g2_nand3_1
X_08997_ _01873_ _01709_ _02654_ VPWR VGND _02743_ sg13g2_or3_1
X_08998_ _02742_ _02743_ _02656_ VPWR VGND _02744_ sg13g2_a21oi_1
X_08999_ _02739_ _02741_ _02744_ VPWR VGND _02745_ sg13g2_a21oi_1
X_09000_ _02677_ _02665_ VPWR VGND _02746_ sg13g2_and2_1
X_09001_ _02745_ _02679_ _02737_ _02746_ VPWR VGND 
+ _02747_
+ sg13g2_a22oi_1
X_09002_ _02044_ _02598_ _02638_ VPWR VGND _02748_ sg13g2_a21oi_1
X_09003_ _02343_ _02599_ VPWR VGND _02749_ sg13g2_xnor2_1
X_09004_ _02748_ _02749_ VPWR VGND _02750_ sg13g2_xnor2_1
X_09005_ _02049_ _02659_ _02738_ _02747_ _02750_ VPWR 
+ VGND
+ _02751_ sg13g2_a221oi_1
X_09006_ _01881_ _01890_ VPWR VGND _02752_ sg13g2_nor2_1
X_09007_ _02278_ _02752_ _02750_ VPWR VGND _02753_ sg13g2_mux2_1
X_09008_ _02049_ _02659_ _02738_ _02747_ _02069_ VPWR 
+ VGND
+ _02754_ sg13g2_a221oi_1
X_09009_ _02652_ _02751_ _02753_ _02754_ VPWR VGND 
+ _02755_
+ sg13g2_or4_1
X_09010_ _02639_ _02640_ VPWR VGND _02756_ sg13g2_nor2_1
X_09011_ _02756_ _02646_ VPWR VGND _02757_ sg13g2_xnor2_1
X_09012_ _02086_ _02757_ VPWR VGND _02758_ sg13g2_nand2_1
X_09013_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2097_o[0]\ VPWR VGND _02759_ sg13g2_buf_1
X_09014_ _02759_ _01902_ VPWR VGND _02760_ sg13g2_and2_1
X_09015_ _02755_ _02758_ _02760_ VPWR VGND _02761_ sg13g2_nand3_1
X_09016_ _02641_ _02756_ _02089_ VPWR VGND _02762_ sg13g2_o21ai_1
X_09017_ _02641_ _02756_ VPWR VGND _02763_ sg13g2_nand2_1
X_09018_ _02762_ _02763_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2099_o\ VPWR VGND _02764_ sg13g2_a21oi_1
X_09019_ _02592_ _02096_ _02764_ _02760_ VPWR VGND 
+ _02765_
+ sg13g2_a22oi_1
X_09020_ _02761_ _02765_ VPWR VGND _00440_ sg13g2_nand2_1
X_09021_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2097_o[1]\ VPWR VGND _02766_ sg13g2_buf_1
X_09022_ _02766_ VPWR VGND _02767_ sg13g2_inv_1
X_09023_ _02767_ _01106_ VPWR VGND _02768_ sg13g2_nor2_1
X_09024_ _02755_ _02758_ _02768_ VPWR VGND _02769_ sg13g2_nand3_1
X_09025_ _02596_ _02096_ _02764_ _02768_ VPWR VGND 
+ _02770_
+ sg13g2_a22oi_1
X_09026_ _02769_ _02770_ VPWR VGND _00441_ sg13g2_nand2_1
X_09027_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2070_o[1]\ VPWR VGND _02771_ sg13g2_buf_1
X_09028_ _02771_ _01244_ VPWR VGND _02772_ sg13g2_nand2_1
X_09029_ \atbs_core_0.comp_lower_sync\ _00864_ _00867_ _00880_ VPWR VGND 
+ _02773_
+ sg13g2_nor4_1
X_09030_ _01244_ _02773_ VPWR VGND _02774_ sg13g2_nand2_1
X_09031_ _01900_ _02772_ _02774_ VPWR VGND _00442_ sg13g2_o21ai_1
X_09032_ _02759_ _02590_ VPWR VGND _02775_ sg13g2_nand2_1
X_09033_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2100_o[0]\ VPWR VGND _02776_ sg13g2_buf_1
X_09034_ _02776_ _02593_ VPWR VGND _02777_ sg13g2_nand2_1
X_09035_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[17]\ VPWR VGND _02778_ sg13g2_inv_1
X_09036_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[14]\ VPWR VGND _02779_ sg13g2_buf_1
X_09037_ _02779_ VPWR VGND _02780_ sg13g2_inv_1
X_09038_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[15]\ VPWR VGND _02781_ sg13g2_buf_1
X_09039_ _01658_ _02781_ VPWR VGND _02782_ sg13g2_nor2_1
X_09040_ _02780_ _02782_ VPWR VGND _02783_ sg13g2_nor2_1
X_09041_ _01675_ _02782_ VPWR VGND _02784_ sg13g2_nor2_1
X_09042_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[12]\ VPWR VGND _02785_ sg13g2_buf_1
X_09043_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[11]\ VPWR VGND _02786_ sg13g2_inv_1
X_09044_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[10]\ VPWR VGND _02787_ sg13g2_buf_1
X_09045_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[8]\ VPWR VGND _02788_ sg13g2_buf_1
X_09046_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[6]\ VPWR VGND _02789_ sg13g2_buf_1
X_09047_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[7]\ VPWR VGND _02790_ sg13g2_buf_1
X_09048_ _01608_ _02789_ _02790_ VPWR VGND _02791_ sg13g2_a21o_1
X_09049_ _02791_ VPWR VGND _02792_ sg13g2_buf_1
X_09050_ _01608_ _02790_ _02789_ VPWR VGND _02793_ sg13g2_and3_1
X_09051_ _02793_ VPWR VGND _02794_ sg13g2_buf_1
X_09052_ _01605_ _02788_ _02792_ _01614_ _02794_ VPWR 
+ VGND
+ _02795_ sg13g2_a221oi_1
X_09053_ _02795_ VPWR VGND _02796_ sg13g2_buf_1
X_09054_ _01619_ _02788_ VPWR VGND _02797_ sg13g2_nor2_1
X_09055_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[9]\ VPWR VGND _02798_ sg13g2_inv_1
X_09056_ _02796_ _02797_ _02798_ VPWR VGND _02799_ sg13g2_o21ai_1
X_09057_ _02798_ _02796_ _02797_ VPWR VGND _02800_ sg13g2_nor3_1
X_09058_ _01604_ _02799_ _02800_ VPWR VGND _02801_ sg13g2_a21o_1
X_09059_ _02801_ VPWR VGND _02802_ sg13g2_buf_1
X_09060_ _02787_ _02802_ VPWR VGND _02803_ sg13g2_nand2_1
X_09061_ _02787_ _02802_ _01648_ VPWR VGND _02804_ sg13g2_o21ai_1
X_09062_ _02786_ _02803_ _02804_ VPWR VGND _02805_ sg13g2_nand3_1
X_09063_ _02803_ _02804_ _02786_ VPWR VGND _02806_ sg13g2_a21oi_1
X_09064_ _01662_ _02785_ _02805_ _01666_ _02806_ VPWR 
+ VGND
+ _02807_ sg13g2_a221oi_1
X_09065_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[13]\ VPWR VGND _02808_ sg13g2_buf_1
X_09066_ _01711_ _02808_ VPWR VGND _02809_ sg13g2_or2_1
X_09067_ _01662_ _02785_ _02809_ VPWR VGND _02810_ sg13g2_o21ai_1
X_09068_ _01712_ _02808_ VPWR VGND _02811_ sg13g2_nand2_1
X_09069_ _02807_ _02810_ _02811_ VPWR VGND _02812_ sg13g2_o21ai_1
X_09070_ _02812_ VPWR VGND _02813_ sg13g2_buf_1
X_09071_ _02783_ _02784_ _02813_ VPWR VGND _02814_ sg13g2_o21ai_1
X_09072_ _02334_ _02780_ _02782_ VPWR VGND _02815_ sg13g2_nor3_1
X_09073_ _01595_ _02781_ _02815_ VPWR VGND _02816_ sg13g2_a21oi_1
X_09074_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[16]\ VPWR VGND _02817_ sg13g2_inv_1
X_09075_ _02814_ _02816_ _02817_ VPWR VGND _02818_ sg13g2_a21oi_1
X_09076_ _02817_ _02814_ _02816_ VPWR VGND _02819_ sg13g2_nand3_1
X_09077_ _02064_ _02818_ _02819_ VPWR VGND _02820_ sg13g2_o21ai_1
X_09078_ _02778_ _02820_ VPWR VGND _02821_ sg13g2_xnor2_1
X_09079_ _01697_ _02821_ VPWR VGND _02822_ sg13g2_xnor2_1
X_09080_ _02086_ _02822_ VPWR VGND _02823_ sg13g2_nand2_1
X_09081_ _02785_ VPWR VGND _02824_ sg13g2_inv_1
X_09082_ _01717_ _02805_ _02806_ VPWR VGND _02825_ sg13g2_a21oi_1
X_09083_ _02824_ _02825_ VPWR VGND _02826_ sg13g2_nand2_1
X_09084_ _02824_ _02825_ _02419_ VPWR VGND _02827_ sg13g2_o21ai_1
X_09085_ _02826_ _02827_ VPWR VGND _02828_ sg13g2_nand2_1
X_09086_ _01946_ _02808_ VPWR VGND _02829_ sg13g2_xor2_1
X_09087_ _02828_ _02829_ VPWR VGND _02830_ sg13g2_xnor2_1
X_09088_ _02575_ _02830_ VPWR VGND _02831_ sg13g2_nand2_1
X_09089_ _01729_ _02787_ VPWR VGND _02832_ sg13g2_xor2_1
X_09090_ _02802_ _02832_ VPWR VGND _02833_ sg13g2_xnor2_1
X_09091_ _01727_ _02833_ VPWR VGND _02834_ sg13g2_nand2_1
X_09092_ _02796_ _02797_ VPWR VGND _02835_ sg13g2_nor2_1
X_09093_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[9]\ VPWR VGND _02836_ sg13g2_xor2_1
X_09094_ _02835_ _02836_ VPWR VGND _02837_ sg13g2_xor2_1
X_09095_ _01959_ _02792_ _02794_ VPWR VGND _02838_ sg13g2_a21oi_1
X_09096_ _01990_ _02788_ VPWR VGND _02839_ sg13g2_xnor2_1
X_09097_ _02838_ _02839_ VPWR VGND _02840_ sg13g2_xnor2_1
X_09098_ _01814_ _02840_ VPWR VGND _02841_ sg13g2_nand2_1
X_09099_ _01812_ _02837_ _02841_ VPWR VGND _02842_ sg13g2_o21ai_1
X_09100_ _02789_ _01774_ VPWR VGND _02843_ sg13g2_xnor2_1
X_09101_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ _02843_ VPWR VGND _02844_ sg13g2_nor2b_1
X_09102_ _01810_ _02843_ VPWR VGND _02845_ sg13g2_and2_1
X_09103_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[193]\ VPWR VGND _02846_ sg13g2_inv_1
X_09104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ VPWR VGND _02847_ sg13g2_inv_1
X_09105_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[191]\ VPWR VGND _02848_ sg13g2_inv_1
X_09106_ _01970_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ VPWR VGND _02849_ sg13g2_nand2b_1
X_09107_ _02848_ _02849_ VPWR VGND _02850_ sg13g2_nand2_1
X_09108_ _02848_ _02849_ VPWR VGND _02851_ sg13g2_nor2_1
X_09109_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ _02850_ _01797_ _02851_ VPWR 
+ VGND
+ _02852_ sg13g2_a221oi_1
X_09110_ _01802_ _02846_ _02847_ _02382_ _02852_ VPWR 
+ VGND
+ _02853_ sg13g2_a221oi_1
X_09111_ _01964_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ VPWR VGND _02854_ sg13g2_nand2_1
X_09112_ _01803_ _02846_ _02854_ VPWR VGND _02855_ sg13g2_o21ai_1
X_09113_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ _01784_ VPWR VGND _02856_ sg13g2_nand2b_1
X_09114_ _02853_ _02855_ _02856_ VPWR VGND _02857_ sg13g2_o21ai_1
X_09115_ _02844_ _02845_ _02857_ VPWR VGND _02858_ sg13g2_o21ai_1
X_09116_ _01957_ _02789_ VPWR VGND _02859_ sg13g2_xnor2_1
X_09117_ _01980_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ VPWR VGND _02860_ sg13g2_nor2_1
X_09118_ _01767_ _02790_ VPWR VGND _02861_ sg13g2_xor2_1
X_09119_ _01957_ _02789_ _02861_ VPWR VGND _02862_ sg13g2_a21o_1
X_09120_ _01819_ _02789_ _02861_ VPWR VGND _02863_ sg13g2_nand3_1
X_09121_ _02862_ _02863_ _01956_ VPWR VGND _02864_ sg13g2_a21oi_1
X_09122_ _01827_ _02859_ _02843_ _02860_ _02864_ VPWR 
+ VGND
+ _02865_ sg13g2_a221oi_1
X_09123_ _02788_ _01756_ VPWR VGND _02866_ sg13g2_xnor2_1
X_09124_ _01840_ _02794_ _02792_ VPWR VGND _02867_ sg13g2_o21ai_1
X_09125_ _01780_ _02867_ VPWR VGND _02868_ sg13g2_nand2_1
X_09126_ _01956_ _02792_ _02868_ VPWR VGND _02869_ sg13g2_o21ai_1
X_09127_ _01819_ _01840_ _02789_ VPWR VGND _02870_ sg13g2_nand3_1
X_09128_ _01959_ _02790_ _02870_ VPWR VGND _02871_ sg13g2_nand3_1
X_09129_ _02863_ _02871_ _02866_ VPWR VGND _02872_ sg13g2_a21oi_1
X_09130_ _02866_ _02869_ _02872_ VPWR VGND _02873_ sg13g2_a21oi_1
X_09131_ _02858_ _02865_ _02873_ VPWR VGND _02874_ sg13g2_a21oi_1
X_09132_ _02787_ _01750_ VPWR VGND _02875_ sg13g2_xnor2_1
X_09133_ _01739_ _02800_ _02799_ VPWR VGND _02876_ sg13g2_o21ai_1
X_09134_ _01739_ _02799_ VPWR VGND _02877_ sg13g2_nor2_1
X_09135_ _01744_ _02876_ _02877_ VPWR VGND _02878_ sg13g2_a21oi_1
X_09136_ _01744_ _02798_ VPWR VGND _02879_ sg13g2_nor2_1
X_09137_ _01739_ _02835_ VPWR VGND _02880_ sg13g2_nand2_1
X_09138_ _02879_ _02880_ _02836_ _02835_ _02875_ VPWR 
+ VGND
+ _02881_ sg13g2_a221oi_1
X_09139_ _02875_ _02878_ _02881_ VPWR VGND _02882_ sg13g2_a21oi_1
X_09140_ _02842_ _02874_ _02882_ VPWR VGND _02883_ sg13g2_o21ai_1
X_09141_ _02834_ _02883_ _02731_ VPWR VGND _02884_ sg13g2_a21oi_1
X_09142_ _02803_ _02804_ VPWR VGND _02885_ sg13g2_nand2_1
X_09143_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[11]\ VPWR VGND _02886_ sg13g2_xor2_1
X_09144_ _02885_ _02886_ VPWR VGND _02887_ sg13g2_xnor2_1
X_09145_ _02731_ _02834_ _02883_ VPWR VGND _02888_ sg13g2_nand3_1
X_09146_ _02884_ _02887_ _02888_ VPWR VGND _02889_ sg13g2_o21ai_1
X_09147_ _01719_ _02785_ VPWR VGND _02890_ sg13g2_xnor2_1
X_09148_ _02825_ _02890_ VPWR VGND _02891_ sg13g2_xnor2_1
X_09149_ _02571_ _02891_ VPWR VGND _02892_ sg13g2_xnor2_1
X_09150_ _01954_ _02891_ VPWR VGND _02893_ sg13g2_nand2_1
X_09151_ _02889_ _02892_ _02893_ VPWR VGND _02894_ sg13g2_o21ai_1
X_09152_ _02575_ _02830_ VPWR VGND _02895_ sg13g2_nor2_1
X_09153_ _02831_ _02894_ _02895_ VPWR VGND _02896_ sg13g2_a21oi_1
X_09154_ _01873_ _02779_ VPWR VGND _02897_ sg13g2_xor2_1
X_09155_ _02813_ _02897_ VPWR VGND _02898_ sg13g2_xnor2_1
X_09156_ _02428_ _02898_ VPWR VGND _02899_ sg13g2_nand2_1
X_09157_ _02049_ _02898_ VPWR VGND _02900_ sg13g2_nand2_1
X_09158_ _02896_ _02899_ _02900_ VPWR VGND _02901_ sg13g2_o21ai_1
X_09159_ _02428_ _02898_ _02896_ VPWR VGND _02902_ sg13g2_nor3_1
X_09160_ _01873_ _02813_ _02779_ VPWR VGND _02903_ sg13g2_a21o_1
X_09161_ _02050_ _02813_ _02903_ VPWR VGND _02904_ sg13g2_o21ai_1
X_09162_ _02044_ _02781_ VPWR VGND _02905_ sg13g2_xor2_1
X_09163_ _02904_ _02905_ VPWR VGND _02906_ sg13g2_xnor2_1
X_09164_ _02814_ _02816_ VPWR VGND _02907_ sg13g2_nand2_1
X_09165_ _02064_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[16]\ VPWR VGND _02908_ sg13g2_xnor2_1
X_09166_ _02907_ _02908_ VPWR VGND _02909_ sg13g2_xnor2_1
X_09167_ _02909_ _01890_ VPWR VGND _02910_ sg13g2_nand2b_1
X_09168_ _02276_ _02906_ _02910_ VPWR VGND _02911_ sg13g2_o21ai_1
X_09169_ _02901_ _02902_ _02911_ VPWR VGND _02912_ sg13g2_nor3_1
X_09170_ _02278_ _02909_ VPWR VGND _02913_ sg13g2_xnor2_1
X_09171_ _02910_ _02906_ VPWR VGND _02914_ sg13g2_and2_1
X_09172_ _02088_ _01689_ VPWR VGND _02915_ sg13g2_xnor2_1
X_09173_ _02915_ _02821_ VPWR VGND _02916_ sg13g2_xnor2_1
X_09174_ _02910_ _02913_ _02914_ _02276_ _02916_ VPWR 
+ VGND
+ _02917_ sg13g2_a221oi_1
X_09175_ _02912_ _02917_ VPWR VGND _02918_ sg13g2_nand2b_1
X_09176_ _02778_ _02820_ _01697_ VPWR VGND _02919_ sg13g2_a21oi_1
X_09177_ _02778_ _02820_ VPWR VGND _02920_ sg13g2_nor2_1
X_09178_ _02919_ _02920_ VPWR VGND _02921_ sg13g2_nor2_1
X_09179_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2102_o\ _02921_ _01902_ VPWR VGND _02922_ sg13g2_o21ai_1
X_09180_ _02823_ _02918_ _02922_ VPWR VGND _02923_ sg13g2_a21oi_1
X_09181_ _02775_ _02777_ _02923_ VPWR VGND _00443_ sg13g2_a21oi_1
X_09182_ _01106_ VPWR VGND _02924_ sg13g2_buf_1
X_09183_ _02766_ _02924_ VPWR VGND _02925_ sg13g2_nand2_1
X_09184_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2100_o[1]\ VPWR VGND _02926_ sg13g2_buf_1
X_09185_ _02926_ _01903_ VPWR VGND _02927_ sg13g2_nand2_1
X_09186_ _02925_ _02927_ _02923_ VPWR VGND _00444_ sg13g2_a21oi_1
X_09187_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[17]\ VPWR VGND _02928_ sg13g2_buf_1
X_09188_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[16]\ VPWR VGND _02929_ sg13g2_buf_1
X_09189_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[15]\ VPWR VGND _02930_ sg13g2_buf_1
X_09190_ _01595_ _02930_ VPWR VGND _02931_ sg13g2_and2_1
X_09191_ _02931_ VPWR VGND _02932_ sg13g2_buf_1
X_09192_ _01658_ _02930_ VPWR VGND _02933_ sg13g2_or2_1
X_09193_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[11]\ VPWR VGND _02934_ sg13g2_inv_1
X_09194_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[10]\ VPWR VGND _02935_ sg13g2_buf_1
X_09195_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[9]\ VPWR VGND _02936_ sg13g2_buf_1
X_09196_ _02936_ VPWR VGND _02937_ sg13g2_inv_1
X_09197_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[8]\ VPWR VGND _02938_ sg13g2_buf_1
X_09198_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[6]\ VPWR VGND _02939_ sg13g2_buf_1
X_09199_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[7]\ VPWR VGND _02940_ sg13g2_buf_1
X_09200_ _01608_ _02939_ _02940_ VPWR VGND _02941_ sg13g2_a21oi_1
X_09201_ _01608_ _02940_ _02939_ VPWR VGND _02942_ sg13g2_nand3_1
X_09202_ _01779_ _02941_ _02942_ VPWR VGND _02943_ sg13g2_o21ai_1
X_09203_ _02943_ VPWR VGND _02944_ sg13g2_buf_1
X_09204_ _02938_ _02944_ VPWR VGND _02945_ sg13g2_nand2_1
X_09205_ _02938_ _02944_ _01606_ VPWR VGND _02946_ sg13g2_o21ai_1
X_09206_ _02937_ _02945_ _02946_ VPWR VGND _02947_ sg13g2_nand3_1
X_09207_ _02945_ _02946_ _02937_ VPWR VGND _02948_ sg13g2_a21oi_1
X_09208_ _01603_ _02947_ _02948_ VPWR VGND _02949_ sg13g2_a21o_1
X_09209_ _02949_ VPWR VGND _02950_ sg13g2_buf_1
X_09210_ _02935_ _02950_ VPWR VGND _02951_ sg13g2_nand2_1
X_09211_ _02935_ _02950_ _01648_ VPWR VGND _02952_ sg13g2_o21ai_1
X_09212_ _02934_ _02951_ _02952_ VPWR VGND _02953_ sg13g2_nand3_1
X_09213_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[12]\ VPWR VGND _02954_ sg13g2_buf_1
X_09214_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[13]\ VPWR VGND _02955_ sg13g2_buf_1
X_09215_ _01599_ _02955_ VPWR VGND _02956_ sg13g2_nand2_1
X_09216_ _02954_ _02956_ VPWR VGND _02957_ sg13g2_nand2b_1
X_09217_ _01915_ _02956_ VPWR VGND _02958_ sg13g2_nand2_1
X_09218_ _02951_ _02952_ _02934_ VPWR VGND _02959_ sg13g2_a21oi_1
X_09219_ _01666_ _02953_ _02957_ _02958_ _02959_ VPWR 
+ VGND
+ _02960_ sg13g2_a221oi_1
X_09220_ _02960_ VPWR VGND _02961_ sg13g2_buf_1
X_09221_ _01661_ _02954_ VPWR VGND _02962_ sg13g2_or2_1
X_09222_ _02962_ _02956_ VPWR VGND _02963_ sg13g2_nand2b_1
X_09223_ _01711_ _02955_ _02963_ VPWR VGND _02964_ sg13g2_o21ai_1
X_09224_ _02964_ VPWR VGND _02965_ sg13g2_buf_1
X_09225_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[14]\ VPWR VGND _02966_ sg13g2_buf_1
X_09226_ _02966_ VPWR VGND _02967_ sg13g2_inv_1
X_09227_ _02961_ _02965_ _02967_ VPWR VGND _02968_ sg13g2_o21ai_1
X_09228_ _02961_ _02965_ _01675_ VPWR VGND _02969_ sg13g2_o21ai_1
X_09229_ _01675_ _02967_ VPWR VGND _02970_ sg13g2_nand2_1
X_09230_ _02933_ _02968_ _02969_ _02970_ VPWR VGND 
+ _02971_
+ sg13g2_and4_1
X_09231_ _02971_ VPWR VGND _02972_ sg13g2_buf_1
X_09232_ _02929_ _02932_ _02972_ VPWR VGND _02973_ sg13g2_nor3_1
X_09233_ _02932_ _02972_ _02929_ VPWR VGND _02974_ sg13g2_o21ai_1
X_09234_ _02491_ _02973_ _02974_ VPWR VGND _02975_ sg13g2_o21ai_1
X_09235_ _02975_ VPWR VGND _02976_ sg13g2_buf_2
X_09236_ _02928_ _02976_ VPWR VGND _02977_ sg13g2_nand2_1
X_09237_ _01697_ _02977_ _01894_ VPWR VGND _02978_ sg13g2_o21ai_1
X_09238_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2105_o\ VPWR VGND _02979_ sg13g2_buf_1
X_09239_ _02928_ _02976_ _02077_ VPWR VGND _02980_ sg13g2_o21ai_1
X_09240_ _01697_ _02977_ _02978_ _02979_ _02980_ VPWR 
+ VGND
+ _02981_ sg13g2_a221oi_1
X_09241_ _02932_ _02972_ VPWR VGND _02982_ sg13g2_or2_1
X_09242_ _02073_ _02929_ VPWR VGND _02983_ sg13g2_nor2_1
X_09243_ _02928_ _02979_ VPWR VGND _02984_ sg13g2_nand2_1
X_09244_ _02088_ _02983_ _02984_ VPWR VGND _02985_ sg13g2_nor3_1
X_09245_ _02073_ _02928_ _02929_ VPWR VGND _02986_ sg13g2_nand3_1
X_09246_ _02928_ _02976_ _02986_ VPWR VGND _02987_ sg13g2_o21ai_1
X_09247_ _02987_ _01697_ VPWR VGND _02988_ sg13g2_nand2b_1
X_09248_ _02928_ _02976_ VPWR VGND _02989_ sg13g2_xnor2_1
X_09249_ _02088_ _02989_ VPWR VGND _02990_ sg13g2_nand2_1
X_09250_ _02982_ _02985_ _02988_ _02990_ _02077_ VPWR 
+ VGND
+ _02991_ sg13g2_a221oi_1
X_09251_ _02088_ _02928_ VPWR VGND _02992_ sg13g2_xor2_1
X_09252_ _02976_ _02992_ VPWR VGND _02993_ sg13g2_xnor2_1
X_09253_ _02064_ _02929_ VPWR VGND _02994_ sg13g2_xor2_1
X_09254_ _02982_ _02994_ VPWR VGND _02995_ sg13g2_xnor2_1
X_09255_ _01658_ _02930_ VPWR VGND _02996_ sg13g2_xor2_1
X_09256_ _02966_ _02996_ VPWR VGND _02997_ sg13g2_and2_1
X_09257_ _01872_ _02996_ VPWR VGND _02998_ sg13g2_and2_1
X_09258_ _02961_ _02965_ VPWR VGND _02999_ sg13g2_nor2_1
X_09259_ _02997_ _02998_ _02999_ VPWR VGND _03000_ sg13g2_o21ai_1
X_09260_ _02966_ _02999_ _02996_ VPWR VGND _03001_ sg13g2_or3_1
X_09261_ _01872_ _02999_ _02996_ VPWR VGND _03002_ sg13g2_or3_1
X_09262_ _03000_ _03001_ _03002_ VPWR VGND _03003_ sg13g2_nand3_1
X_09263_ _01873_ _02966_ _02996_ VPWR VGND _03004_ sg13g2_nand3_1
X_09264_ _02970_ _02996_ _03004_ VPWR VGND _03005_ sg13g2_o21ai_1
X_09265_ _03003_ _03005_ _01887_ VPWR VGND _03006_ sg13g2_o21ai_1
X_09266_ _01871_ _02966_ VPWR VGND _03007_ sg13g2_xnor2_1
X_09267_ _02961_ _02965_ _03007_ VPWR VGND _03008_ sg13g2_o21ai_1
X_09268_ _02961_ _02965_ _03007_ VPWR VGND _03009_ sg13g2_or3_1
X_09269_ _03008_ _03009_ _01703_ VPWR VGND _03010_ sg13g2_a21oi_1
X_09270_ _01667_ _02953_ _02959_ VPWR VGND _03011_ sg13g2_a21o_1
X_09271_ _01951_ _02954_ VPWR VGND _03012_ sg13g2_and2_1
X_09272_ _03011_ _02962_ _03012_ VPWR VGND _03013_ sg13g2_a21oi_1
X_09273_ _01946_ _02955_ VPWR VGND _03014_ sg13g2_xnor2_1
X_09274_ _03013_ _03014_ VPWR VGND _03015_ sg13g2_xnor2_1
X_09275_ _01913_ _03015_ VPWR VGND _03016_ sg13g2_nor2_1
X_09276_ _01719_ _02954_ VPWR VGND _03017_ sg13g2_xor2_1
X_09277_ _03011_ _03017_ VPWR VGND _03018_ sg13g2_xnor2_1
X_09278_ _01856_ _03018_ VPWR VGND _03019_ sg13g2_xnor2_1
X_09279_ _02935_ _01750_ VPWR VGND _03020_ sg13g2_xor2_1
X_09280_ _02945_ _02946_ VPWR VGND _03021_ sg13g2_nand2_1
X_09281_ _01735_ _02936_ VPWR VGND _03022_ sg13g2_xor2_1
X_09282_ _01736_ _02936_ VPWR VGND _03023_ sg13g2_nand2_1
X_09283_ _01738_ _03021_ _03023_ VPWR VGND _03024_ sg13g2_a21oi_1
X_09284_ _03021_ _03022_ _03024_ VPWR VGND _03025_ sg13g2_a21oi_1
X_09285_ _02936_ _03021_ VPWR VGND _03026_ sg13g2_nor2_1
X_09286_ _01738_ _02948_ _02947_ VPWR VGND _03027_ sg13g2_o21ai_1
X_09287_ _02687_ _03026_ _03027_ _01744_ _03020_ VPWR 
+ VGND
+ _03028_ sg13g2_a221oi_1
X_09288_ _03020_ _03025_ _03028_ VPWR VGND _03029_ sg13g2_a21oi_1
X_09289_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ VPWR VGND _03030_ sg13g2_buf_1
X_09290_ _03030_ _02234_ _01834_ VPWR VGND _03031_ sg13g2_o21ai_1
X_09291_ _01764_ _02939_ VPWR VGND _03032_ sg13g2_xnor2_1
X_09292_ _03031_ _03032_ VPWR VGND _03033_ sg13g2_and2_1
X_09293_ _03030_ _02238_ _03032_ VPWR VGND _03034_ sg13g2_nor3_1
X_09294_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ VPWR VGND _03035_ sg13g2_nor2b_1
X_09295_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _03035_ VPWR VGND _03036_ sg13g2_nand2_1
X_09296_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _03035_ _01796_ VPWR VGND _03037_ sg13g2_o21ai_1
X_09297_ _01965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ VPWR VGND _03038_ sg13g2_nand2_1
X_09298_ _03036_ _03037_ _03038_ VPWR VGND _03039_ sg13g2_nand3_1
X_09299_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ VPWR VGND _03040_ sg13g2_inv_1
X_09300_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ _01783_ VPWR VGND _03041_ sg13g2_nand2b_1
X_09301_ _02221_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _03041_ VPWR VGND _03042_ sg13g2_o21ai_1
X_09302_ _01787_ _03040_ _03042_ VPWR VGND _03043_ sg13g2_a21oi_1
X_09303_ _01783_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ VPWR VGND _03044_ sg13g2_nor2b_1
X_09304_ _01801_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ VPWR VGND _03045_ sg13g2_nor2b_1
X_09305_ _03044_ _03045_ _03041_ VPWR VGND _03046_ sg13g2_o21ai_1
X_09306_ _01809_ _03030_ VPWR VGND _03047_ sg13g2_xnor2_1
X_09307_ _02939_ _01773_ VPWR VGND _03048_ sg13g2_xnor2_1
X_09308_ _03046_ _03047_ _03048_ VPWR VGND _03049_ sg13g2_nand3_1
X_09309_ _03039_ _03043_ _03049_ VPWR VGND _03050_ sg13g2_a21oi_1
X_09310_ _03033_ _03034_ _03050_ VPWR VGND _03051_ sg13g2_nor3_1
X_09311_ _01819_ _02939_ VPWR VGND _03052_ sg13g2_nand2_1
X_09312_ _01759_ _02940_ VPWR VGND _03053_ sg13g2_xor2_1
X_09313_ _03052_ _03053_ VPWR VGND _03054_ sg13g2_xnor2_1
X_09314_ _01956_ _03051_ _03054_ VPWR VGND _03055_ sg13g2_o21ai_1
X_09315_ _02938_ _02944_ VPWR VGND _03056_ sg13g2_xnor2_1
X_09316_ _01756_ _03056_ VPWR VGND _03057_ sg13g2_xnor2_1
X_09317_ _01956_ _03051_ _03057_ VPWR VGND _03058_ sg13g2_a21oi_1
X_09318_ _03021_ _03022_ VPWR VGND _03059_ sg13g2_xor2_1
X_09319_ _01990_ _03056_ VPWR VGND _03060_ sg13g2_xor2_1
X_09320_ _01814_ _03060_ VPWR VGND _03061_ sg13g2_nand2_1
X_09321_ _01739_ _03059_ _03061_ VPWR VGND _03062_ sg13g2_o21ai_1
X_09322_ _03055_ _03058_ _03062_ VPWR VGND _03063_ sg13g2_a21o_1
X_09323_ _01729_ _02935_ VPWR VGND _03064_ sg13g2_xor2_1
X_09324_ _02950_ _03064_ VPWR VGND _03065_ sg13g2_xnor2_1
X_09325_ _03029_ _03063_ _03065_ _01727_ VPWR VGND 
+ _03066_
+ sg13g2_a22oi_1
X_09326_ _02731_ _03066_ VPWR VGND _03067_ sg13g2_nand2_1
X_09327_ _02951_ _02952_ VPWR VGND _03068_ sg13g2_nand2_1
X_09328_ _01717_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[11]\ VPWR VGND _03069_ sg13g2_xnor2_1
X_09329_ _03068_ _03069_ VPWR VGND _03070_ sg13g2_xnor2_1
X_09330_ _02731_ _03066_ _03070_ VPWR VGND _03071_ sg13g2_o21ai_1
X_09331_ _03067_ _03071_ VPWR VGND _03072_ sg13g2_and2_1
X_09332_ _01722_ _03018_ _03019_ _03072_ _01913_ VPWR 
+ VGND
+ _03073_ sg13g2_a221oi_1
X_09333_ _01722_ _03018_ _03019_ _03072_ _03015_ VPWR 
+ VGND
+ _03074_ sg13g2_a221oi_1
X_09334_ _03008_ _03009_ VPWR VGND _03075_ sg13g2_nand2_1
X_09335_ _02428_ _03075_ VPWR VGND _03076_ sg13g2_xor2_1
X_09336_ _03016_ _03073_ _03074_ _03076_ VPWR VGND 
+ _03077_
+ sg13g2_nor4_1
X_09337_ _01887_ _03003_ _03005_ VPWR VGND _03078_ sg13g2_or3_1
X_09338_ _03010_ _03077_ _03078_ VPWR VGND _03079_ sg13g2_o21ai_1
X_09339_ _01881_ _02995_ VPWR VGND _03080_ sg13g2_or2_1
X_09340_ _02278_ _02995_ VPWR VGND _03081_ sg13g2_nand2_1
X_09341_ _03006_ _03079_ _03080_ _03081_ VPWR VGND 
+ _03082_
+ sg13g2_a22oi_1
X_09342_ _02086_ _02993_ _02995_ _02069_ _03082_ VPWR 
+ VGND
+ _03083_ sg13g2_a221oi_1
X_09343_ _02088_ _02928_ _02976_ VPWR VGND _03084_ sg13g2_nor3_1
X_09344_ _01691_ _03084_ VPWR VGND _03085_ sg13g2_and2_1
X_09345_ _02077_ _02979_ _03084_ VPWR VGND _03086_ sg13g2_nor3_1
X_09346_ _01105_ _03085_ _03086_ VPWR VGND _03087_ sg13g2_or3_1
X_09347_ _02981_ _02991_ _03083_ _03087_ VPWR VGND 
+ _03088_
+ sg13g2_or4_1
X_09348_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2103_o[0]\ VPWR VGND _03089_ sg13g2_buf_1
X_09349_ _03089_ VPWR VGND _03090_ sg13g2_inv_1
X_09350_ _02776_ _02589_ VPWR VGND _03091_ sg13g2_nand2_1
X_09351_ _03090_ _02103_ _03091_ VPWR VGND _03092_ sg13g2_o21ai_1
X_09352_ _03088_ _03092_ VPWR VGND _00445_ sg13g2_and2_1
X_09353_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2103_o[1]\ VPWR VGND _03093_ sg13g2_buf_1
X_09354_ _03093_ VPWR VGND _03094_ sg13g2_inv_1
X_09355_ _02926_ _02589_ VPWR VGND _03095_ sg13g2_nand2_1
X_09356_ _03094_ _02103_ _03095_ VPWR VGND _03096_ sg13g2_o21ai_1
X_09357_ _03088_ _03096_ VPWR VGND _00446_ sg13g2_and2_1
X_09358_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2106_o[0]\ VPWR VGND _03097_ sg13g2_buf_1
X_09359_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[6]\ VPWR VGND _03098_ sg13g2_buf_1
X_09360_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[7]\ VPWR VGND _03099_ sg13g2_buf_1
X_09361_ _01609_ _03098_ _03099_ VPWR VGND _03100_ sg13g2_a21o_1
X_09362_ _01763_ _03099_ _03098_ VPWR VGND _03101_ sg13g2_and3_1
X_09363_ _01959_ _03100_ _03101_ VPWR VGND _03102_ sg13g2_a21oi_1
X_09364_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[8]\ VPWR VGND _03103_ sg13g2_buf_1
X_09365_ _01990_ _03103_ VPWR VGND _03104_ sg13g2_xnor2_1
X_09366_ _03102_ _03104_ VPWR VGND _03105_ sg13g2_xnor2_1
X_09367_ _01767_ _03099_ VPWR VGND _03106_ sg13g2_xnor2_1
X_09368_ _01761_ _01834_ VPWR VGND _03107_ sg13g2_nand2_1
X_09369_ _01957_ _03098_ _03107_ VPWR VGND _03108_ sg13g2_nand3_1
X_09370_ _01840_ _01837_ VPWR VGND _03109_ sg13g2_nor2_1
X_09371_ _03098_ _03109_ VPWR VGND _03110_ sg13g2_nand2b_1
X_09372_ _03106_ _03108_ _03110_ VPWR VGND _03111_ sg13g2_o21ai_1
X_09373_ _03098_ _01826_ VPWR VGND _03112_ sg13g2_nand2b_1
X_09374_ _01841_ _03112_ _01957_ VPWR VGND _03113_ sg13g2_a21oi_1
X_09375_ _01983_ _03098_ _01841_ VPWR VGND _03114_ sg13g2_a21oi_1
X_09376_ _03113_ _03114_ _03106_ VPWR VGND _03115_ sg13g2_o21ai_1
X_09377_ _03111_ _03115_ VPWR VGND _03116_ sg13g2_nor2b_1
X_09378_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[233]\ VPWR VGND _03117_ sg13g2_inv_1
X_09379_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ VPWR VGND _03118_ sg13g2_inv_1
X_09380_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ VPWR VGND _03119_ sg13g2_inv_1
X_09381_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[229]\ VPWR VGND _03120_ sg13g2_inv_1
X_09382_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ VPWR VGND _03121_ sg13g2_nand2b_1
X_09383_ _03120_ _03121_ VPWR VGND _03122_ sg13g2_nand2_1
X_09384_ _03120_ _03121_ VPWR VGND _03123_ sg13g2_nor2_1
X_09385_ _01965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ _03122_ _01797_ _03123_ VPWR 
+ VGND
+ _03124_ sg13g2_a221oi_1
X_09386_ _01802_ _03118_ _03119_ _01788_ _03124_ VPWR 
+ VGND
+ _03125_ sg13g2_a221oi_1
X_09387_ _01963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ VPWR VGND _03126_ sg13g2_nand2_1
X_09388_ _01802_ _03118_ _03126_ VPWR VGND _03127_ sg13g2_o21ai_1
X_09389_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ _01783_ VPWR VGND _03128_ sg13g2_nand2b_1
X_09390_ _03125_ _03127_ _03128_ VPWR VGND _03129_ sg13g2_o21ai_1
X_09391_ _03117_ _03129_ _01810_ VPWR VGND _03130_ sg13g2_o21ai_1
X_09392_ _03117_ _03129_ VPWR VGND _03131_ sg13g2_nand2_1
X_09393_ _01832_ _01771_ VPWR VGND _03132_ sg13g2_nand2_1
X_09394_ _03106_ _03132_ VPWR VGND _03133_ sg13g2_xnor2_1
X_09395_ _03098_ _01774_ VPWR VGND _03134_ sg13g2_xnor2_1
X_09396_ _02548_ _03133_ _03134_ VPWR VGND _03135_ sg13g2_o21ai_1
X_09397_ _03130_ _03131_ _03135_ VPWR VGND _03136_ sg13g2_a21o_1
X_09398_ _03105_ _01989_ VPWR VGND _03137_ sg13g2_nand2b_1
X_09399_ _01754_ _03105_ VPWR VGND _03138_ sg13g2_nand2_1
X_09400_ _03116_ _03136_ _03137_ _03138_ VPWR VGND 
+ _03139_
+ sg13g2_a22oi_1
X_09401_ _01998_ _03105_ _03139_ VPWR VGND _03140_ sg13g2_a21oi_1
X_09402_ _01606_ _03103_ _03100_ _01614_ _03101_ VPWR 
+ VGND
+ _03141_ sg13g2_a221oi_1
X_09403_ _01606_ _03103_ VPWR VGND _03142_ sg13g2_nor2_1
X_09404_ _03141_ _03142_ VPWR VGND _03143_ sg13g2_nor2_1
X_09405_ _01740_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[9]\ VPWR VGND _03144_ sg13g2_xor2_1
X_09406_ _03143_ _03144_ VPWR VGND _03145_ sg13g2_xnor2_1
X_09407_ _03145_ VPWR VGND _03146_ sg13g2_inv_1
X_09408_ _02001_ _03140_ _03146_ VPWR VGND _03147_ sg13g2_o21ai_1
X_09409_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[9]\ VPWR VGND _03148_ sg13g2_inv_1
X_09410_ _03141_ _03142_ _03148_ VPWR VGND _03149_ sg13g2_o21ai_1
X_09411_ _03148_ _03141_ _03142_ VPWR VGND _03150_ sg13g2_nor3_1
X_09412_ _01604_ _03149_ _03150_ VPWR VGND _03151_ sg13g2_a21o_1
X_09413_ _03151_ VPWR VGND _03152_ sg13g2_buf_1
X_09414_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[10]\ VPWR VGND _03153_ sg13g2_buf_1
X_09415_ _01730_ _03153_ VPWR VGND _03154_ sg13g2_xor2_1
X_09416_ _03152_ _03154_ VPWR VGND _03155_ sg13g2_xnor2_1
X_09417_ _02197_ _03155_ VPWR VGND _03156_ sg13g2_or2_1
X_09418_ _02001_ _03140_ _03156_ VPWR VGND _03157_ sg13g2_a21oi_1
X_09419_ _03147_ _03157_ _02015_ VPWR VGND _03158_ sg13g2_a21oi_1
X_09420_ _03153_ _03152_ VPWR VGND _03159_ sg13g2_nand2_1
X_09421_ _03153_ _03152_ _01648_ VPWR VGND _03160_ sg13g2_o21ai_1
X_09422_ _03159_ _03160_ VPWR VGND _03161_ sg13g2_nand2_1
X_09423_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[11]\ VPWR VGND _03162_ sg13g2_xor2_1
X_09424_ _03161_ _03162_ VPWR VGND _03163_ sg13g2_xnor2_1
X_09425_ _03147_ _03157_ _03163_ VPWR VGND _03164_ sg13g2_a21oi_1
X_09426_ _02197_ _03145_ VPWR VGND _03165_ sg13g2_nand2_1
X_09427_ _02197_ _02687_ VPWR VGND _03166_ sg13g2_nand2_1
X_09428_ _03165_ _03166_ _03140_ VPWR VGND _03167_ sg13g2_a21oi_1
X_09429_ _03146_ _03166_ _01728_ VPWR VGND _03168_ sg13g2_o21ai_1
X_09430_ _03167_ _03168_ _03155_ VPWR VGND _03169_ sg13g2_o21ai_1
X_09431_ _03158_ _03164_ _03169_ VPWR VGND _03170_ sg13g2_o21ai_1
X_09432_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[12]\ VPWR VGND _03171_ sg13g2_buf_1
X_09433_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[11]\ VPWR VGND _03172_ sg13g2_inv_1
X_09434_ _03172_ _03159_ _03160_ VPWR VGND _03173_ sg13g2_nand3_1
X_09435_ _03159_ _03160_ _03172_ VPWR VGND _03174_ sg13g2_a21oi_1
X_09436_ _01666_ _03173_ _03174_ VPWR VGND _03175_ sg13g2_a21o_1
X_09437_ _03175_ VPWR VGND _03176_ sg13g2_buf_1
X_09438_ _03171_ _03176_ VPWR VGND _03177_ sg13g2_xnor2_1
X_09439_ _01858_ _03177_ VPWR VGND _03178_ sg13g2_xnor2_1
X_09440_ _02015_ _03163_ VPWR VGND _03179_ sg13g2_nor2_1
X_09441_ _03178_ _03179_ VPWR VGND _03180_ sg13g2_nor2_1
X_09442_ _03171_ _03176_ VPWR VGND _03181_ sg13g2_nand2_1
X_09443_ _03171_ _03176_ _01662_ VPWR VGND _03182_ sg13g2_o21ai_1
X_09444_ _03181_ _03182_ VPWR VGND _03183_ sg13g2_nand2_1
X_09445_ _01947_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[13]\ VPWR VGND _03184_ sg13g2_xnor2_1
X_09446_ _03183_ _03184_ VPWR VGND _03185_ sg13g2_xnor2_1
X_09447_ _02419_ _03177_ VPWR VGND _03186_ sg13g2_xnor2_1
X_09448_ _01954_ _03186_ VPWR VGND _03187_ sg13g2_nand2_1
X_09449_ _03185_ _03187_ VPWR VGND _03188_ sg13g2_nand2_1
X_09450_ _02575_ _03187_ VPWR VGND _03189_ sg13g2_nand2_1
X_09451_ _03170_ _03180_ _03188_ _03189_ VPWR VGND 
+ _03190_
+ sg13g2_a22oi_1
X_09452_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[15]\ VPWR VGND _03191_ sg13g2_buf_1
X_09453_ _01876_ _03191_ VPWR VGND _03192_ sg13g2_xnor2_1
X_09454_ _03192_ VPWR VGND _03193_ sg13g2_buf_1
X_09455_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[14]\ VPWR VGND _03194_ sg13g2_buf_1
X_09456_ _01709_ _03194_ VPWR VGND _03195_ sg13g2_or2_1
X_09457_ _02428_ _03194_ _03193_ VPWR VGND _03196_ sg13g2_nand3_1
X_09458_ _03193_ _03195_ _03196_ VPWR VGND _03197_ sg13g2_o21ai_1
X_09459_ _01709_ _03194_ _03193_ VPWR VGND _03198_ sg13g2_a21o_1
X_09460_ _01887_ _03198_ _02334_ VPWR VGND _03199_ sg13g2_o21ai_1
X_09461_ _02036_ _03193_ _03195_ VPWR VGND _03200_ sg13g2_nand3_1
X_09462_ _02050_ _03200_ VPWR VGND _03201_ sg13g2_nand2_1
X_09463_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[13]\ VPWR VGND _03202_ sg13g2_inv_1
X_09464_ _01912_ _03202_ VPWR VGND _03203_ sg13g2_nor2_1
X_09465_ _01912_ _03202_ _03181_ _03182_ VPWR VGND 
+ _03204_
+ sg13g2_a22oi_1
X_09466_ _03203_ _03204_ VPWR VGND _03205_ sg13g2_nor2_1
X_09467_ _01709_ _03194_ VPWR VGND _03206_ sg13g2_xnor2_1
X_09468_ _03205_ _03206_ VPWR VGND _03207_ sg13g2_xnor2_1
X_09469_ _03199_ _03201_ _03207_ VPWR VGND _03208_ sg13g2_mux2_1
X_09470_ _02037_ _03197_ _03185_ _02575_ _03208_ VPWR 
+ VGND
+ _03209_ sg13g2_a221oi_1
X_09471_ _03190_ _03209_ VPWR VGND _03210_ sg13g2_nand2b_1
X_09472_ _01912_ _03202_ VPWR VGND _03211_ sg13g2_nand2_1
X_09473_ _01658_ _03191_ VPWR VGND _03212_ sg13g2_nand2_1
X_09474_ _01912_ _03202_ _03212_ VPWR VGND _03213_ sg13g2_o21ai_1
X_09475_ _01871_ _03194_ _03211_ _03183_ _03213_ VPWR 
+ VGND
+ _03214_ sg13g2_a221oi_1
X_09476_ _01706_ _03194_ VPWR VGND _03215_ sg13g2_nor2_1
X_09477_ _01876_ _03191_ VPWR VGND _03216_ sg13g2_nor2_1
X_09478_ _03212_ _03215_ _03216_ VPWR VGND _03217_ sg13g2_a21oi_1
X_09479_ _03214_ _03217_ VPWR VGND _03218_ sg13g2_nand2b_1
X_09480_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[16]\ VPWR VGND _03219_ sg13g2_buf_1
X_09481_ _02064_ _03219_ VPWR VGND _03220_ sg13g2_xnor2_1
X_09482_ _03218_ _03220_ VPWR VGND _03221_ sg13g2_xnor2_1
X_09483_ _01873_ _03194_ VPWR VGND _03222_ sg13g2_xor2_1
X_09484_ _03205_ _03222_ _02048_ VPWR VGND _03223_ sg13g2_o21ai_1
X_09485_ _02050_ _03194_ VPWR VGND _03224_ sg13g2_nand2_1
X_09486_ _02048_ _03205_ _03224_ VPWR VGND _03225_ sg13g2_a21oi_1
X_09487_ _03203_ _03204_ _01703_ VPWR VGND _03226_ sg13g2_o21ai_1
X_09488_ _01887_ _03226_ _03215_ VPWR VGND _03227_ sg13g2_a21oi_1
X_09489_ _03225_ _03227_ VPWR VGND _03228_ sg13g2_or2_1
X_09490_ _01886_ _02047_ VPWR VGND _03229_ sg13g2_nand2_1
X_09491_ _03229_ _03203_ _03204_ VPWR VGND _03230_ sg13g2_nor3_1
X_09492_ _03230_ _03215_ VPWR VGND _03231_ sg13g2_nand2b_1
X_09493_ _03205_ _03222_ VPWR VGND _03232_ sg13g2_nand2_1
X_09494_ _03231_ _03232_ _03193_ VPWR VGND _03233_ sg13g2_a21oi_1
X_09495_ _02037_ _03223_ _03228_ _03193_ _03233_ VPWR 
+ VGND
+ _03234_ sg13g2_a221oi_1
X_09496_ _02069_ _03221_ _03234_ VPWR VGND _03235_ sg13g2_a21oi_1
X_09497_ _03210_ _03235_ VPWR VGND _03236_ sg13g2_nand2_1
X_09498_ _01681_ _03219_ VPWR VGND _03237_ sg13g2_nand2_1
X_09499_ _02064_ _03219_ VPWR VGND _03238_ sg13g2_nor2_1
X_09500_ _03218_ _03237_ _03238_ VPWR VGND _03239_ sg13g2_a21o_1
X_09501_ _03239_ VPWR VGND _03240_ sg13g2_buf_1
X_09502_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2108_o\ VPWR VGND _03241_ sg13g2_inv_1
X_09503_ _03241_ _00949_ _03218_ _03237_ _03238_ VPWR 
+ VGND
+ _03242_ sg13g2_a221oi_1
X_09504_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[17]\ VPWR VGND _03243_ sg13g2_buf_1
X_09505_ _03240_ _03242_ _03243_ VPWR VGND _03244_ sg13g2_mux2_1
X_09506_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2108_o\ _01105_ VPWR VGND _03245_ sg13g2_nor2_1
X_09507_ _02289_ _03245_ _02290_ VPWR VGND _03246_ sg13g2_o21ai_1
X_09508_ _03243_ _03240_ VPWR VGND _03247_ sg13g2_xnor2_1
X_09509_ _02292_ _03244_ _03246_ _03247_ VPWR VGND 
+ _03248_
+ sg13g2_a22oi_1
X_09510_ _02278_ _03221_ VPWR VGND _03249_ sg13g2_xnor2_1
X_09511_ _01890_ _03221_ _03249_ VPWR VGND _03250_ sg13g2_a21oi_1
X_09512_ _03248_ _03250_ VPWR VGND _03251_ sg13g2_nor2_1
X_09513_ _01895_ _03241_ VPWR VGND _03252_ sg13g2_nor2_1
X_09514_ _03243_ VPWR VGND _03253_ sg13g2_inv_1
X_09515_ _03253_ _03240_ VPWR VGND _03254_ sg13g2_or2_1
X_09516_ _02089_ _03247_ VPWR VGND _03255_ sg13g2_nand2_1
X_09517_ _02089_ _03254_ _03255_ VPWR VGND _03256_ sg13g2_o21ai_1
X_09518_ _02088_ _01894_ _03243_ VPWR VGND _03257_ sg13g2_nor3_1
X_09519_ _03240_ _03257_ _01106_ VPWR VGND _03258_ sg13g2_a21o_1
X_09520_ _03236_ _03251_ _03252_ _03256_ _03258_ VPWR 
+ VGND
+ _03259_ sg13g2_a221oi_1
X_09521_ _03090_ _01903_ VPWR VGND _03260_ sg13g2_nor2_1
X_09522_ _03097_ _03259_ _03260_ VPWR VGND _00447_ sg13g2_a21o_1
X_09523_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2106_o[1]\ VPWR VGND _03261_ sg13g2_buf_1
X_09524_ _03094_ _01903_ VPWR VGND _03262_ sg13g2_nor2_1
X_09525_ _03261_ _03259_ _03262_ VPWR VGND _00448_ sg13g2_a21o_1
X_09526_ _03097_ VPWR VGND _03263_ sg13g2_inv_1
X_09527_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2109_o[0]\ VPWR VGND _03264_ sg13g2_buf_1
X_09528_ _03264_ _01902_ VPWR VGND _03265_ sg13g2_nand2_1
X_09529_ _03263_ _02108_ _03265_ VPWR VGND _03266_ sg13g2_o21ai_1
X_09530_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[16]\ VPWR VGND _03267_ sg13g2_buf_1
X_09531_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[15]\ VPWR VGND _03268_ sg13g2_buf_1
X_09532_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[14]\ VPWR VGND _03269_ sg13g2_buf_1
X_09533_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[12]\ VPWR VGND _03270_ sg13g2_buf_1
X_09534_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[11]\ VPWR VGND _03271_ sg13g2_inv_1
X_09535_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[13]\ VPWR VGND _03272_ sg13g2_buf_1
X_09536_ _01599_ _03272_ VPWR VGND _03273_ sg13g2_nand2_1
X_09537_ _01916_ _03271_ _03273_ VPWR VGND _03274_ sg13g2_o21ai_1
X_09538_ _03270_ _03274_ VPWR VGND _03275_ sg13g2_or2_1
X_09539_ _03274_ _01915_ VPWR VGND _03276_ sg13g2_nand2b_1
X_09540_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[10]\ VPWR VGND _03277_ sg13g2_buf_1
X_09541_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[9]\ VPWR VGND _03278_ sg13g2_inv_1
X_09542_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[8]\ VPWR VGND _03279_ sg13g2_buf_1
X_09543_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[6]\ VPWR VGND _03280_ sg13g2_buf_1
X_09544_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[7]\ VPWR VGND _03281_ sg13g2_buf_1
X_09545_ _01763_ _03280_ _03281_ VPWR VGND _03282_ sg13g2_a21oi_1
X_09546_ _01763_ _03281_ _03280_ VPWR VGND _03283_ sg13g2_nand3_1
X_09547_ _01780_ _03282_ _03283_ VPWR VGND _03284_ sg13g2_o21ai_1
X_09548_ _03279_ _03284_ VPWR VGND _03285_ sg13g2_nand2_1
X_09549_ _03279_ _03284_ _01619_ VPWR VGND _03286_ sg13g2_o21ai_1
X_09550_ _03278_ _03285_ _03286_ VPWR VGND _03287_ sg13g2_nand3_1
X_09551_ _03285_ _03286_ _03278_ VPWR VGND _03288_ sg13g2_a21oi_1
X_09552_ _01604_ _03287_ _03288_ VPWR VGND _03289_ sg13g2_a21o_1
X_09553_ _03289_ VPWR VGND _03290_ sg13g2_buf_1
X_09554_ _03277_ _03290_ VPWR VGND _03291_ sg13g2_nand2_1
X_09555_ _03277_ _03290_ _01729_ VPWR VGND _03292_ sg13g2_o21ai_1
X_09556_ _02018_ _03271_ _03291_ _03292_ VPWR VGND 
+ _03293_
+ sg13g2_a22oi_1
X_09557_ _03275_ _03276_ _03293_ VPWR VGND _03294_ sg13g2_a21o_1
X_09558_ _01661_ _03270_ VPWR VGND _03295_ sg13g2_nor2_1
X_09559_ _01711_ _03272_ VPWR VGND _03296_ sg13g2_nor2_1
X_09560_ _03273_ _03295_ _03296_ VPWR VGND _03297_ sg13g2_a21oi_1
X_09561_ _03269_ _03294_ _03297_ VPWR VGND _03298_ sg13g2_nand3_1
X_09562_ _03294_ _03297_ _03269_ VPWR VGND _03299_ sg13g2_a21oi_1
X_09563_ _02334_ _03298_ _03299_ VPWR VGND _03300_ sg13g2_a21oi_1
X_09564_ _03268_ _03300_ _01876_ VPWR VGND _03301_ sg13g2_a21o_1
X_09565_ _03301_ VPWR VGND _03302_ sg13g2_buf_1
X_09566_ _03268_ _03300_ VPWR VGND _03303_ sg13g2_or2_1
X_09567_ _03303_ VPWR VGND _03304_ sg13g2_buf_1
X_09568_ _03267_ _03302_ _03304_ VPWR VGND _03305_ sg13g2_nand3_1
X_09569_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[17]\ VPWR VGND _03306_ sg13g2_buf_1
X_09570_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2111_o\ VPWR VGND _03307_ sg13g2_inv_1
X_09571_ _03306_ _03307_ VPWR VGND _03308_ sg13g2_nand2_1
X_09572_ _01686_ _03307_ VPWR VGND _03309_ sg13g2_nand2_1
X_09573_ _03302_ _03304_ _03267_ VPWR VGND _03310_ sg13g2_a21oi_1
X_09574_ _02491_ _03305_ _03308_ _03309_ _03310_ VPWR 
+ VGND
+ _03311_ sg13g2_a221oi_1
X_09575_ _01686_ _03306_ VPWR VGND _03312_ sg13g2_nand2_1
X_09576_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2111_o\ _03312_ _00949_ VPWR VGND _03313_ sg13g2_o21ai_1
X_09577_ _03311_ _03313_ VPWR VGND _03314_ sg13g2_or2_1
X_09578_ _02491_ _03305_ _03310_ VPWR VGND _03315_ sg13g2_a21oi_1
X_09579_ _01686_ _03306_ VPWR VGND _03316_ sg13g2_xnor2_1
X_09580_ _03315_ _03316_ VPWR VGND _03317_ sg13g2_xnor2_1
X_09581_ _02077_ _03314_ _03317_ VPWR VGND _03318_ sg13g2_nor3_1
X_09582_ _03311_ _03313_ VPWR VGND _03319_ sg13g2_nor2_1
X_09583_ _02077_ _03319_ _03317_ VPWR VGND _03320_ sg13g2_and3_1
X_09584_ _02018_ _03271_ VPWR VGND _03321_ sg13g2_nor2_1
X_09585_ _03270_ _03321_ _03293_ VPWR VGND _03322_ sg13g2_nor3_1
X_09586_ _03321_ _03293_ _03270_ VPWR VGND _03323_ sg13g2_o21ai_1
X_09587_ _03322_ _03323_ VPWR VGND _03324_ sg13g2_nor2b_1
X_09588_ _01951_ _03324_ VPWR VGND _03325_ sg13g2_xnor2_1
X_09589_ _02419_ _03322_ _03323_ VPWR VGND _03326_ sg13g2_o21ai_1
X_09590_ _01946_ _03272_ VPWR VGND _03327_ sg13g2_xnor2_1
X_09591_ _03326_ _03327_ VPWR VGND _03328_ sg13g2_xnor2_1
X_09592_ _02575_ _03328_ VPWR VGND _03329_ sg13g2_nor2_1
X_09593_ _01954_ _03325_ _03329_ VPWR VGND _03330_ sg13g2_a21oi_1
X_09594_ _03291_ _03292_ VPWR VGND _03331_ sg13g2_nand2_1
X_09595_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[11]\ VPWR VGND _03332_ sg13g2_xnor2_1
X_09596_ _03331_ _03332_ VPWR VGND _03333_ sg13g2_xnor2_1
X_09597_ _01990_ _03279_ VPWR VGND _03334_ sg13g2_xnor2_1
X_09598_ _03284_ _03334_ VPWR VGND _03335_ sg13g2_xnor2_1
X_09599_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[252]\ VPWR VGND _03336_ sg13g2_inv_1
X_09600_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ VPWR VGND _03337_ sg13g2_inv_1
X_09601_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ VPWR VGND _03338_ sg13g2_inv_1
X_09602_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[248]\ VPWR VGND _03339_ sg13g2_inv_1
X_09603_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ VPWR VGND _03340_ sg13g2_nand2b_1
X_09604_ _03339_ _03340_ VPWR VGND _03341_ sg13g2_nand2_1
X_09605_ _03339_ _03340_ VPWR VGND _03342_ sg13g2_nor2_1
X_09606_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ _03341_ _01797_ _03342_ VPWR 
+ VGND
+ _03343_ sg13g2_a221oi_1
X_09607_ _01802_ _03337_ _03338_ _02382_ _03343_ VPWR 
+ VGND
+ _03344_ sg13g2_a221oi_1
X_09608_ _01963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ VPWR VGND _03345_ sg13g2_nand2_1
X_09609_ _01802_ _03337_ _03345_ VPWR VGND _03346_ sg13g2_o21ai_1
X_09610_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ _01783_ VPWR VGND _03347_ sg13g2_nand2b_1
X_09611_ _03344_ _03346_ _03347_ VPWR VGND _03348_ sg13g2_o21ai_1
X_09612_ _01810_ _03336_ _03348_ VPWR VGND _03349_ sg13g2_a21o_1
X_09613_ _03280_ _01774_ VPWR VGND _03350_ sg13g2_xor2_1
X_09614_ _01980_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[252]\ _03350_ VPWR VGND _03351_ sg13g2_a21oi_1
X_09615_ _01758_ _03281_ VPWR VGND _03352_ sg13g2_xnor2_1
X_09616_ _02548_ _03352_ VPWR VGND _03353_ sg13g2_nand2_1
X_09617_ _01957_ _03280_ VPWR VGND _03354_ sg13g2_xor2_1
X_09618_ _01956_ _01983_ _03353_ _03354_ VPWR VGND 
+ _03355_
+ sg13g2_a22oi_1
X_09619_ _01819_ _03280_ VPWR VGND _03356_ sg13g2_nand2_1
X_09620_ _01957_ _03356_ _03352_ VPWR VGND _03357_ sg13g2_mux2_1
X_09621_ _01827_ _03357_ VPWR VGND _03358_ sg13g2_or2_1
X_09622_ _03349_ _03351_ _03355_ _03358_ VPWR VGND 
+ _03359_
+ sg13g2_a22oi_1
X_09623_ _02548_ _03280_ _03352_ VPWR VGND _03360_ sg13g2_nor3_1
X_09624_ _02548_ _03357_ VPWR VGND _03361_ sg13g2_nor2_1
X_09625_ _03360_ _03361_ VPWR VGND _03362_ sg13g2_or2_1
X_09626_ _01754_ _03359_ _03362_ VPWR VGND _03363_ sg13g2_or3_1
X_09627_ _01998_ _03335_ VPWR VGND _03364_ sg13g2_nor2_1
X_09628_ _01989_ _03359_ _03362_ VPWR VGND _03365_ sg13g2_or3_1
X_09629_ _03277_ _03290_ VPWR VGND _03366_ sg13g2_xnor2_1
X_09630_ _01750_ _03366_ VPWR VGND _03367_ sg13g2_xor2_1
X_09631_ _03285_ _03286_ VPWR VGND _03368_ sg13g2_nand2_1
X_09632_ _01740_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[9]\ VPWR VGND _03369_ sg13g2_xor2_1
X_09633_ _03368_ _03369_ VPWR VGND _03370_ sg13g2_xnor2_1
X_09634_ _03367_ _03370_ VPWR VGND _03371_ sg13g2_nand2_1
X_09635_ _03335_ _03363_ _03364_ _03365_ _03371_ VPWR 
+ VGND
+ _03372_ sg13g2_a221oi_1
X_09636_ _02687_ _03367_ VPWR VGND _03373_ sg13g2_nand2_1
X_09637_ _03335_ _03363_ _03364_ _03365_ _03373_ VPWR 
+ VGND
+ _03374_ sg13g2_a221oi_1
X_09638_ _01628_ _03366_ VPWR VGND _03375_ sg13g2_xnor2_1
X_09639_ _02250_ _03375_ VPWR VGND _03376_ sg13g2_nand2_1
X_09640_ _02001_ _03371_ _03376_ VPWR VGND _03377_ sg13g2_o21ai_1
X_09641_ _03372_ _03374_ _03377_ VPWR VGND _03378_ sg13g2_nor3_1
X_09642_ _03333_ _03378_ VPWR VGND _03379_ sg13g2_nand2_1
X_09643_ _03333_ _03378_ _02731_ VPWR VGND _03380_ sg13g2_o21ai_1
X_09644_ _03379_ _03380_ VPWR VGND _03381_ sg13g2_nand2_1
X_09645_ _03330_ _03381_ VPWR VGND _03382_ sg13g2_nand2_1
X_09646_ _01858_ _03324_ VPWR VGND _03383_ sg13g2_xor2_1
X_09647_ _03294_ _03297_ VPWR VGND _03384_ sg13g2_nand2_1
X_09648_ _01873_ _03269_ VPWR VGND _03385_ sg13g2_xnor2_1
X_09649_ _03384_ _03385_ VPWR VGND _03386_ sg13g2_xnor2_1
X_09650_ _02428_ _03386_ VPWR VGND _03387_ sg13g2_xor2_1
X_09651_ _02575_ _03328_ _03330_ _03383_ _03387_ VPWR 
+ VGND
+ _03388_ sg13g2_a221oi_1
X_09652_ _02044_ _03268_ VPWR VGND _03389_ sg13g2_xnor2_1
X_09653_ _03300_ _03389_ VPWR VGND _03390_ sg13g2_xnor2_1
X_09654_ _02049_ _03386_ VPWR VGND _03391_ sg13g2_nand2_1
X_09655_ _03390_ _03391_ VPWR VGND _03392_ sg13g2_nand2_1
X_09656_ _02276_ _03391_ VPWR VGND _03393_ sg13g2_nand2_1
X_09657_ _03268_ _03300_ _02044_ VPWR VGND _03394_ sg13g2_a21oi_1
X_09658_ _03268_ _03300_ VPWR VGND _03395_ sg13g2_nor2_1
X_09659_ _01890_ VPWR VGND _03396_ sg13g2_inv_1
X_09660_ _01682_ _03267_ VPWR VGND _03397_ sg13g2_xor2_1
X_09661_ _03396_ _03397_ VPWR VGND _03398_ sg13g2_nor2_1
X_09662_ _03394_ _03395_ _03398_ VPWR VGND _03399_ sg13g2_o21ai_1
X_09663_ _01890_ _03302_ _03304_ _03397_ VPWR VGND 
+ _03400_
+ sg13g2_nand4_1
X_09664_ _03399_ _03400_ VPWR VGND _03401_ sg13g2_nand2_1
X_09665_ _03382_ _03388_ _03392_ _03393_ _03401_ VPWR 
+ VGND
+ _03402_ sg13g2_a221oi_1
X_09666_ _01881_ _03397_ VPWR VGND _03403_ sg13g2_nand2_1
X_09667_ _01682_ _03267_ VPWR VGND _03404_ sg13g2_xnor2_1
X_09668_ _01881_ _03404_ VPWR VGND _03405_ sg13g2_nand2b_1
X_09669_ _03302_ _03304_ _03403_ _03405_ VPWR VGND 
+ _03406_
+ sg13g2_a22oi_1
X_09670_ _01881_ _03394_ _03395_ _03404_ VPWR VGND 
+ _03407_
+ sg13g2_nor4_1
X_09671_ _01881_ _03302_ _03304_ _03404_ VPWR VGND 
+ _03408_
+ sg13g2_and4_1
X_09672_ _03406_ _03407_ _03408_ VPWR VGND _03409_ sg13g2_nor3_1
X_09673_ _02276_ _03390_ VPWR VGND _03410_ sg13g2_nand2_1
X_09674_ _03409_ _03410_ _03401_ VPWR VGND _03411_ sg13g2_a21oi_1
X_09675_ _03402_ _03411_ VPWR VGND _03412_ sg13g2_nor2_1
X_09676_ _03318_ _03320_ _03412_ VPWR VGND _03413_ sg13g2_o21ai_1
X_09677_ _01895_ _03314_ _03317_ VPWR VGND _03414_ sg13g2_or3_1
X_09678_ _03266_ _03413_ _03414_ VPWR VGND _00449_ sg13g2_and3_1
X_09679_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2109_o[1]\ VPWR VGND _03415_ sg13g2_buf_1
X_09680_ _03415_ VPWR VGND _03416_ sg13g2_inv_1
X_09681_ _03261_ _02589_ VPWR VGND _03417_ sg13g2_nand2_1
X_09682_ _03416_ _01107_ _03417_ VPWR VGND _03418_ sg13g2_o21ai_1
X_09683_ _03413_ _03414_ _03418_ VPWR VGND _00450_ sg13g2_and3_1
X_09684_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[12]\ VPWR VGND _03419_ sg13g2_buf_1
X_09685_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[11]\ VPWR VGND _03420_ sg13g2_inv_1
X_09686_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[10]\ VPWR VGND _03421_ sg13g2_buf_1
X_09687_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[9]\ VPWR VGND _03422_ sg13g2_inv_1
X_09688_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[8]\ VPWR VGND _03423_ sg13g2_buf_1
X_09689_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[6]\ VPWR VGND _03424_ sg13g2_buf_1
X_09690_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[7]\ VPWR VGND _03425_ sg13g2_buf_1
X_09691_ _01608_ _03424_ _03425_ VPWR VGND _03426_ sg13g2_a21o_1
X_09692_ _01608_ _03425_ _03424_ VPWR VGND _03427_ sg13g2_and3_1
X_09693_ _01614_ _03426_ _03427_ VPWR VGND _03428_ sg13g2_a21o_1
X_09694_ _03428_ VPWR VGND _03429_ sg13g2_buf_1
X_09695_ _03423_ _03429_ VPWR VGND _03430_ sg13g2_nand2_1
X_09696_ _03423_ _03429_ _01619_ VPWR VGND _03431_ sg13g2_o21ai_1
X_09697_ _03422_ _03430_ _03431_ VPWR VGND _03432_ sg13g2_nand3_1
X_09698_ _03430_ _03431_ _03422_ VPWR VGND _03433_ sg13g2_a21oi_1
X_09699_ _01604_ _03432_ _03433_ VPWR VGND _03434_ sg13g2_a21o_1
X_09700_ _03434_ VPWR VGND _03435_ sg13g2_buf_1
X_09701_ _01648_ _03421_ _03435_ VPWR VGND _03436_ sg13g2_o21ai_1
X_09702_ _01639_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[11]\ _03421_ _01648_ VPWR VGND 
+ _03437_
+ sg13g2_a22oi_1
X_09703_ _01916_ _03420_ _03436_ _03437_ VPWR VGND 
+ _03438_
+ sg13g2_a22oi_1
X_09704_ _03438_ VPWR VGND _03439_ sg13g2_buf_1
X_09705_ _03419_ _03439_ _01662_ VPWR VGND _03440_ sg13g2_a21oi_1
X_09706_ _03419_ _03439_ VPWR VGND _03441_ sg13g2_nor2_1
X_09707_ _03440_ _03441_ VPWR VGND _03442_ sg13g2_nor2_1
X_09708_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[13]\ VPWR VGND _03443_ sg13g2_buf_1
X_09709_ _01947_ _03443_ VPWR VGND _03444_ sg13g2_xor2_1
X_09710_ _03419_ _03439_ _01951_ VPWR VGND _03445_ sg13g2_a21o_1
X_09711_ _03419_ _03439_ VPWR VGND _03446_ sg13g2_or2_1
X_09712_ _03446_ VPWR VGND _03447_ sg13g2_buf_1
X_09713_ _01711_ _03443_ VPWR VGND _03448_ sg13g2_nand2_1
X_09714_ _03445_ _03447_ _03448_ VPWR VGND _03449_ sg13g2_a21oi_1
X_09715_ _03442_ _03444_ _03449_ VPWR VGND _03450_ sg13g2_a21oi_1
X_09716_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[14]\ VPWR VGND _03451_ sg13g2_buf_1
X_09717_ _03451_ _01908_ VPWR VGND _03452_ sg13g2_xnor2_1
X_09718_ _02029_ _03452_ VPWR VGND _03453_ sg13g2_or2_1
X_09719_ _03419_ _03439_ VPWR VGND _03454_ sg13g2_xnor2_1
X_09720_ _02419_ _03454_ VPWR VGND _03455_ sg13g2_xnor2_1
X_09721_ _02030_ _03452_ VPWR VGND _03456_ sg13g2_and2_1
X_09722_ _03445_ _03447_ _03443_ VPWR VGND _03457_ sg13g2_a21oi_1
X_09723_ _01954_ _03455_ _03456_ _03457_ VPWR VGND 
+ _03458_
+ sg13g2_a22oi_1
X_09724_ _03450_ _03453_ _03458_ VPWR VGND _03459_ sg13g2_o21ai_1
X_09725_ _01730_ _03421_ VPWR VGND _03460_ sg13g2_xor2_1
X_09726_ _03435_ _03460_ VPWR VGND _03461_ sg13g2_xnor2_1
X_09727_ _02197_ _03461_ VPWR VGND _03462_ sg13g2_or2_1
X_09728_ _02197_ _03461_ VPWR VGND _03463_ sg13g2_nand2_1
X_09729_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _01784_ VPWR VGND _03464_ sg13g2_nand2b_1
X_09730_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ VPWR VGND _03465_ sg13g2_inv_1
X_09731_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ VPWR VGND _03466_ sg13g2_inv_1
X_09732_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ VPWR VGND _03467_ sg13g2_inv_1
X_09733_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ VPWR VGND _03468_ sg13g2_nand2b_1
X_09734_ _03467_ _03468_ VPWR VGND _03469_ sg13g2_nand2_1
X_09735_ _03467_ _03468_ VPWR VGND _03470_ sg13g2_nor2_1
X_09736_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ _03469_ _01797_ _03470_ VPWR 
+ VGND
+ _03471_ sg13g2_a221oi_1
X_09737_ _01802_ _03465_ _03466_ _02382_ _03471_ VPWR 
+ VGND
+ _03472_ sg13g2_a221oi_1
X_09738_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _01964_ VPWR VGND 
+ _03473_
+ sg13g2_a22oi_1
X_09739_ _03472_ _03473_ VPWR VGND _03474_ sg13g2_nand2b_1
X_09740_ _03424_ _01774_ VPWR VGND _03475_ sg13g2_xor2_1
X_09741_ _01980_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _03464_ _03474_ _03475_ VPWR 
+ VGND
+ _03476_ sg13g2_a221oi_1
X_09742_ _01980_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _03475_ VPWR VGND _03477_ sg13g2_nor3_1
X_09743_ _01819_ _03424_ VPWR VGND _03478_ sg13g2_xnor2_1
X_09744_ _01832_ _03424_ VPWR VGND _03479_ sg13g2_nand2_1
X_09745_ _01767_ _03425_ VPWR VGND _03480_ sg13g2_xor2_1
X_09746_ _03479_ _03480_ VPWR VGND _03481_ sg13g2_xor2_1
X_09747_ _01827_ _03478_ _03481_ _02213_ VPWR VGND 
+ _03482_
+ sg13g2_a22oi_1
X_09748_ _03477_ _03482_ VPWR VGND _03483_ sg13g2_nand2b_1
X_09749_ _03423_ _01756_ VPWR VGND _03484_ sg13g2_xnor2_1
X_09750_ _01840_ _03427_ _03426_ VPWR VGND _03485_ sg13g2_o21ai_1
X_09751_ _01780_ _03485_ VPWR VGND _03486_ sg13g2_nand2_1
X_09752_ _01841_ _03426_ _03486_ VPWR VGND _03487_ sg13g2_o21ai_1
X_09753_ _03479_ _03480_ VPWR VGND _03488_ sg13g2_nand2b_1
X_09754_ _01819_ _01840_ _03424_ VPWR VGND _03489_ sg13g2_nand3_1
X_09755_ _01959_ _03425_ _03489_ VPWR VGND _03490_ sg13g2_nand3_1
X_09756_ _03488_ _03490_ _03484_ VPWR VGND _03491_ sg13g2_a21oi_1
X_09757_ _03484_ _03487_ _03491_ VPWR VGND _03492_ sg13g2_a21o_1
X_09758_ _03476_ _03483_ _03492_ VPWR VGND _03493_ sg13g2_o21ai_1
X_09759_ _01990_ _03423_ VPWR VGND _03494_ sg13g2_xor2_1
X_09760_ _03429_ _03494_ VPWR VGND _03495_ sg13g2_xnor2_1
X_09761_ _01998_ _03495_ VPWR VGND _03496_ sg13g2_nand2_1
X_09762_ _02001_ _03493_ _03496_ VPWR VGND _03497_ sg13g2_nand3_1
X_09763_ _03430_ _03431_ VPWR VGND _03498_ sg13g2_nand2_1
X_09764_ _01740_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[9]\ VPWR VGND _03499_ sg13g2_xor2_1
X_09765_ _03498_ _03499_ VPWR VGND _03500_ sg13g2_xnor2_1
X_09766_ _03493_ _03496_ _02001_ VPWR VGND _03501_ sg13g2_a21oi_1
X_09767_ _03497_ _03500_ _03501_ VPWR VGND _03502_ sg13g2_a21oi_1
X_09768_ _03462_ _03463_ _03502_ VPWR VGND _03503_ sg13g2_a21oi_1
X_09769_ _01730_ _03435_ VPWR VGND _03504_ sg13g2_nand2_1
X_09770_ _01730_ _03435_ _03421_ VPWR VGND _03505_ sg13g2_o21ai_1
X_09771_ _03504_ _03505_ VPWR VGND _03506_ sg13g2_nand2_1
X_09772_ _01717_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[11]\ VPWR VGND _03507_ sg13g2_xnor2_1
X_09773_ _03506_ _03507_ VPWR VGND _03508_ sg13g2_xnor2_1
X_09774_ _02250_ _03461_ VPWR VGND _03509_ sg13g2_nand2_1
X_09775_ _03508_ _03509_ VPWR VGND _03510_ sg13g2_nand2_1
X_09776_ _03503_ _03510_ _02015_ VPWR VGND _03511_ sg13g2_o21ai_1
X_09777_ _03508_ _03502_ _03462_ VPWR VGND _03512_ sg13g2_nor3_1
X_09778_ _03508_ _03502_ _03463_ VPWR VGND _03513_ sg13g2_nor3_1
X_09779_ _03508_ _03509_ VPWR VGND _03514_ sg13g2_nor2_1
X_09780_ _03512_ _03513_ _03514_ VPWR VGND _03515_ sg13g2_nor3_1
X_09781_ _01858_ _03454_ VPWR VGND _03516_ sg13g2_xnor2_1
X_09782_ _03511_ _03515_ _03516_ VPWR VGND _03517_ sg13g2_a21oi_1
X_09783_ _02029_ _03442_ _03448_ VPWR VGND _03518_ sg13g2_a21oi_1
X_09784_ _03442_ _03444_ _03518_ VPWR VGND _03519_ sg13g2_a21o_1
X_09785_ _03443_ _03445_ _03447_ VPWR VGND _03520_ sg13g2_nand3_1
X_09786_ _01725_ _03520_ _03457_ VPWR VGND _03521_ sg13g2_a21oi_1
X_09787_ _01913_ _03457_ VPWR VGND _03522_ sg13g2_nand2_1
X_09788_ _01947_ _03521_ _03522_ VPWR VGND _03523_ sg13g2_o21ai_1
X_09789_ _03519_ _03523_ _03452_ VPWR VGND _03524_ sg13g2_mux2_1
X_09790_ _03459_ _03517_ _03524_ VPWR VGND _03525_ sg13g2_o21ai_1
X_09791_ _01712_ _03443_ VPWR VGND _03526_ sg13g2_or2_1
X_09792_ _03526_ VPWR VGND _03527_ sg13g2_buf_1
X_09793_ _03440_ _03441_ _03448_ VPWR VGND _03528_ sg13g2_o21ai_1
X_09794_ _03528_ VPWR VGND _03529_ sg13g2_buf_1
X_09795_ _03451_ _03527_ _03529_ VPWR VGND _03530_ sg13g2_nand3_1
X_09796_ _03527_ _03529_ _03451_ VPWR VGND _03531_ sg13g2_a21oi_1
X_09797_ _02334_ _03530_ _03531_ VPWR VGND _03532_ sg13g2_a21o_1
X_09798_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[15]\ VPWR VGND _03533_ sg13g2_buf_1
X_09799_ _02044_ _03533_ VPWR VGND _03534_ sg13g2_xor2_1
X_09800_ _03532_ _03534_ VPWR VGND _03535_ sg13g2_xnor2_1
X_09801_ _01873_ _03451_ VPWR VGND _03536_ sg13g2_xor2_1
X_09802_ _03527_ _03529_ _03536_ VPWR VGND _03537_ sg13g2_a21oi_1
X_09803_ _03527_ _03529_ _03536_ VPWR VGND _03538_ sg13g2_and3_1
X_09804_ _03537_ _03538_ _02048_ VPWR VGND _03539_ sg13g2_o21ai_1
X_09805_ _03535_ _03539_ VPWR VGND _03540_ sg13g2_and2_1
X_09806_ _03525_ _03540_ _02276_ VPWR VGND _03541_ sg13g2_a21oi_1
X_09807_ _03525_ _03539_ _03535_ VPWR VGND _03542_ sg13g2_a21oi_1
X_09808_ _01877_ _03533_ VPWR VGND _03543_ sg13g2_nand2_1
X_09809_ _01876_ _03533_ VPWR VGND _03544_ sg13g2_nor2_1
X_09810_ _03532_ _03543_ _03544_ VPWR VGND _03545_ sg13g2_a21o_1
X_09811_ _03545_ VPWR VGND _03546_ sg13g2_buf_1
X_09812_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[16]\ VPWR VGND _03547_ sg13g2_buf_1
X_09813_ _02073_ _03547_ VPWR VGND _03548_ sg13g2_xnor2_1
X_09814_ _03546_ _03548_ VPWR VGND _03549_ sg13g2_xnor2_1
X_09815_ _02278_ _03549_ VPWR VGND _03550_ sg13g2_xnor2_1
X_09816_ _03541_ _03542_ _03550_ VPWR VGND _03551_ sg13g2_o21ai_1
X_09817_ _02069_ _03549_ VPWR VGND _03552_ sg13g2_nand2_1
X_09818_ _03551_ _03552_ VPWR VGND _03553_ sg13g2_nand2_1
X_09819_ _03264_ _01106_ VPWR VGND _03554_ sg13g2_and2_1
X_09820_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[17]\ VPWR VGND _03555_ sg13g2_buf_1
X_09821_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2446_o\ _01105_ VPWR VGND _03556_ sg13g2_nor2_1
X_09822_ _03556_ VPWR VGND _03557_ sg13g2_buf_1
X_09823_ _03555_ _03547_ _03557_ VPWR VGND _03558_ sg13g2_nand3_1
X_09824_ _01685_ _03547_ _03557_ VPWR VGND _03559_ sg13g2_nand3_1
X_09825_ _03558_ _03559_ _03546_ VPWR VGND _03560_ sg13g2_a21oi_1
X_09826_ _02343_ _03555_ _03557_ VPWR VGND _03561_ sg13g2_nand3_1
X_09827_ _01685_ _02343_ _03557_ VPWR VGND _03562_ sg13g2_nand3_1
X_09828_ _03561_ _03562_ _03546_ VPWR VGND _03563_ sg13g2_a21oi_1
X_09829_ _02073_ _03555_ _03547_ _03557_ VPWR VGND 
+ _03564_
+ sg13g2_nand4_1
X_09830_ _01685_ _02343_ _03547_ _03557_ VPWR VGND 
+ _03565_
+ sg13g2_nand4_1
X_09831_ _01686_ _03555_ _03557_ VPWR VGND _03566_ sg13g2_nand3_1
X_09832_ _03564_ _03565_ _03566_ VPWR VGND _03567_ sg13g2_nand3_1
X_09833_ _03560_ _03563_ _03567_ VPWR VGND _03568_ sg13g2_or3_1
X_09834_ _03568_ VPWR VGND _03569_ sg13g2_buf_1
X_09835_ _03547_ VPWR VGND _03570_ sg13g2_inv_1
X_09836_ _03533_ _03451_ _03547_ VPWR VGND _03571_ sg13g2_or3_1
X_09837_ _03451_ VPWR VGND _03572_ sg13g2_inv_1
X_09838_ _01674_ _03572_ _03570_ VPWR VGND _03573_ sg13g2_nand3_1
X_09839_ _03527_ _03529_ _03571_ _03573_ VPWR VGND 
+ _03574_
+ sg13g2_a22oi_1
X_09840_ _01871_ _03533_ VPWR VGND _03575_ sg13g2_nor2_1
X_09841_ _03570_ _03575_ VPWR VGND _03576_ sg13g2_nand2_1
X_09842_ _01876_ _01871_ VPWR VGND _03577_ sg13g2_nor2_1
X_09843_ _03570_ _03577_ VPWR VGND _03578_ sg13g2_nand2_1
X_09844_ _03527_ _03529_ _03576_ _03578_ VPWR VGND 
+ _03579_
+ sg13g2_a22oi_1
X_09845_ _03451_ _03547_ VPWR VGND _03580_ sg13g2_nor2_1
X_09846_ _03577_ _03575_ _03580_ VPWR VGND _03581_ sg13g2_o21ai_1
X_09847_ _03570_ _03544_ VPWR VGND _03582_ sg13g2_nand2_1
X_09848_ _03581_ _03582_ VPWR VGND _03583_ sg13g2_nand2_1
X_09849_ _03574_ _03579_ _03583_ VPWR VGND _03584_ sg13g2_nor3_1
X_09850_ _02073_ _03584_ VPWR VGND _03585_ sg13g2_nand2_1
X_09851_ _03570_ _03546_ _03585_ VPWR VGND _03586_ sg13g2_o21ai_1
X_09852_ _01685_ _03555_ VPWR VGND _03587_ sg13g2_xor2_1
X_09853_ _03586_ _03587_ VPWR VGND _03588_ sg13g2_xor2_1
X_09854_ _01897_ _03588_ VPWR VGND _03589_ sg13g2_xnor2_1
X_09855_ _03554_ _03569_ _03589_ VPWR VGND _03590_ sg13g2_nor3_1
X_09856_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2934_o\ VPWR VGND _03591_ sg13g2_buf_1
X_09857_ _03570_ _03546_ VPWR VGND _03592_ sg13g2_nor2_1
X_09858_ _02086_ _03587_ VPWR VGND _03593_ sg13g2_and2_1
X_09859_ _01894_ _03584_ _03587_ VPWR VGND _03594_ sg13g2_nor3_1
X_09860_ _03592_ _03593_ _03594_ VPWR VGND _03595_ sg13g2_a21oi_1
X_09861_ _02073_ _01894_ _03587_ VPWR VGND _03596_ sg13g2_nor3_1
X_09862_ _03570_ _03546_ _03596_ VPWR VGND _03597_ sg13g2_o21ai_1
X_09863_ _02073_ _01690_ _03584_ _03587_ VPWR VGND 
+ _03598_
+ sg13g2_nand4_1
X_09864_ _00949_ _03597_ _03598_ VPWR VGND _03599_ sg13g2_and3_1
X_09865_ _03595_ _03599_ _03569_ VPWR VGND _03600_ sg13g2_a21o_1
X_09866_ _03591_ _03600_ _03554_ VPWR VGND _03601_ sg13g2_a21oi_1
X_09867_ _03553_ _03590_ _03601_ VPWR VGND _00451_ sg13g2_a21oi_1
X_09868_ _03416_ _01902_ VPWR VGND _03602_ sg13g2_nor2_1
X_09869_ _03569_ _03589_ _03602_ VPWR VGND _03603_ sg13g2_nor3_1
X_09870_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2931_o\ _03600_ _03602_ VPWR VGND _03604_ sg13g2_a21oi_1
X_09871_ _03553_ _03603_ _03604_ VPWR VGND _00452_ sg13g2_a21oi_1
X_09872_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2073_o[0]\ VPWR VGND _03605_ sg13g2_buf_1
X_09873_ _03605_ VPWR VGND _03606_ sg13g2_inv_1
X_09874_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[16]\ VPWR VGND _03607_ sg13g2_buf_1
X_09875_ _02064_ _03607_ VPWR VGND _03608_ sg13g2_nor2_1
X_09876_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[14]\ VPWR VGND _03609_ sg13g2_buf_1
X_09877_ _01672_ _03609_ VPWR VGND _03610_ sg13g2_and2_1
X_09878_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[12]\ VPWR VGND _03611_ sg13g2_buf_1
X_09879_ _03611_ VPWR VGND _03612_ sg13g2_inv_1
X_09880_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[10]\ VPWR VGND _03613_ sg13g2_buf_1
X_09881_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[8]\ VPWR VGND _03614_ sg13g2_buf_1
X_09882_ _01605_ _03614_ VPWR VGND _03615_ sg13g2_nor2_1
X_09883_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[6]\ VPWR VGND _03616_ sg13g2_buf_2
X_09884_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[7]\ VPWR VGND _03617_ sg13g2_buf_1
X_09885_ _01608_ _03616_ _03617_ VPWR VGND _03618_ sg13g2_a21o_1
X_09886_ _01608_ _03617_ _03616_ VPWR VGND _03619_ sg13g2_and3_1
X_09887_ _01605_ _03614_ _03618_ _01613_ _03619_ VPWR 
+ VGND
+ _03620_ sg13g2_a221oi_1
X_09888_ _03620_ VPWR VGND _03621_ sg13g2_buf_1
X_09889_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[9]\ VPWR VGND _03622_ sg13g2_inv_1
X_09890_ _03615_ _03621_ _03622_ VPWR VGND _03623_ sg13g2_o21ai_1
X_09891_ _03623_ VPWR VGND _03624_ sg13g2_buf_2
X_09892_ _03622_ _03615_ _03621_ VPWR VGND _03625_ sg13g2_nor3_1
X_09893_ _01603_ _03624_ _03625_ VPWR VGND _03626_ sg13g2_a21o_1
X_09894_ _03626_ VPWR VGND _03627_ sg13g2_buf_1
X_09895_ _03613_ _03627_ VPWR VGND _03628_ sg13g2_nand2_1
X_09896_ _03613_ _03627_ _01627_ VPWR VGND _03629_ sg13g2_o21ai_1
X_09897_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[11]\ VPWR VGND _03630_ sg13g2_buf_1
X_09898_ _01639_ _03630_ VPWR VGND _03631_ sg13g2_nor2_1
X_09899_ _03628_ _03629_ _03631_ VPWR VGND _03632_ sg13g2_a21o_1
X_09900_ _01639_ _03630_ VPWR VGND _03633_ sg13g2_nand2_1
X_09901_ _03632_ _03633_ VPWR VGND _03634_ sg13g2_and2_1
X_09902_ _03634_ VPWR VGND _03635_ sg13g2_buf_2
X_09903_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[13]\ VPWR VGND _03636_ sg13g2_buf_1
X_09904_ _03609_ _03636_ VPWR VGND _03637_ sg13g2_nand2_1
X_09905_ _01672_ _03636_ VPWR VGND _03638_ sg13g2_nand2_1
X_09906_ _03630_ VPWR VGND _03639_ sg13g2_inv_1
X_09907_ _01916_ _03639_ _03628_ _03629_ _03612_ VPWR 
+ VGND
+ _03640_ sg13g2_a221oi_1
X_09908_ _01916_ _03612_ _03639_ VPWR VGND _03641_ sg13g2_nor3_1
X_09909_ _01662_ _03640_ _03641_ VPWR VGND _03642_ sg13g2_nor3_1
X_09910_ _03612_ _03635_ _03637_ _03638_ _03642_ VPWR 
+ VGND
+ _03643_ sg13g2_a221oi_1
X_09911_ _01712_ _03609_ VPWR VGND _03644_ sg13g2_nand2_1
X_09912_ _01671_ _01712_ VPWR VGND _03645_ sg13g2_nand2_1
X_09913_ _03612_ _03635_ _03644_ _03645_ _03642_ VPWR 
+ VGND
+ _03646_ sg13g2_a221oi_1
X_09914_ _03636_ VPWR VGND _03647_ sg13g2_inv_1
X_09915_ _03644_ _03645_ _03647_ VPWR VGND _03648_ sg13g2_a21oi_1
X_09916_ _03610_ _03643_ _03646_ _03648_ VPWR VGND 
+ _03649_
+ sg13g2_nor4_1
X_09917_ _01658_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[15]\ VPWR VGND _03650_ sg13g2_nand2_1
X_09918_ _01658_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[15]\ VPWR VGND _03651_ sg13g2_nor2_1
X_09919_ _03649_ _03650_ _03651_ VPWR VGND _03652_ sg13g2_a21o_1
X_09920_ _02064_ _03607_ VPWR VGND _03653_ sg13g2_nand2_1
X_09921_ _03608_ _03652_ _03653_ VPWR VGND _03654_ sg13g2_o21ai_1
X_09922_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[17]\ VPWR VGND _03655_ sg13g2_buf_1
X_09923_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2075_o\ _03655_ VPWR VGND _03656_ sg13g2_nor2b_1
X_09924_ _03655_ _03654_ VPWR VGND _03657_ sg13g2_nor2_1
X_09925_ _01696_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2075_o\ _03657_ VPWR VGND _03658_ sg13g2_nor3_1
X_09926_ _03654_ _03656_ _03658_ VPWR VGND _03659_ sg13g2_a21oi_1
X_09927_ _01686_ _03655_ VPWR VGND _03660_ sg13g2_xor2_1
X_09928_ _03654_ _03660_ VPWR VGND _03661_ sg13g2_xnor2_1
X_09929_ _01661_ _03640_ _03641_ VPWR VGND _03662_ sg13g2_or3_1
X_09930_ _03662_ VPWR VGND _03663_ sg13g2_buf_1
X_09931_ _03612_ _03632_ _03633_ VPWR VGND _03664_ sg13g2_nand3_1
X_09932_ _03664_ VPWR VGND _03665_ sg13g2_buf_1
X_09933_ _03663_ _03665_ VPWR VGND _03666_ sg13g2_and2_1
X_09934_ _03666_ VPWR VGND _03667_ sg13g2_buf_2
X_09935_ _01671_ _03609_ VPWR VGND _03668_ sg13g2_xor2_1
X_09936_ _02047_ _03636_ _03667_ _03668_ VPWR VGND 
+ _03669_
+ sg13g2_and4_1
X_09937_ _01713_ _02047_ _03667_ _03668_ VPWR VGND 
+ _03670_
+ sg13g2_and4_1
X_09938_ _01702_ _03647_ VPWR VGND _03671_ sg13g2_nand2_1
X_09939_ _01600_ _01702_ VPWR VGND _03672_ sg13g2_nand2_1
X_09940_ _03663_ _03665_ _03671_ _03672_ _03668_ VPWR 
+ VGND
+ _03673_ sg13g2_a221oi_1
X_09941_ _01712_ _01703_ VPWR VGND _03674_ sg13g2_nor2_1
X_09942_ _03647_ _03674_ VPWR VGND _03675_ sg13g2_nand2_1
X_09943_ _01713_ _02047_ _03636_ _03668_ VPWR VGND 
+ _03676_
+ sg13g2_nand4_1
X_09944_ _03668_ _03675_ _03676_ VPWR VGND _03677_ sg13g2_o21ai_1
X_09945_ _03669_ _03670_ _03673_ _03677_ VPWR VGND 
+ _03678_
+ sg13g2_nor4_1
X_09946_ _03651_ _03650_ VPWR VGND _03679_ sg13g2_nor2b_1
X_09947_ _03649_ _03678_ _03679_ VPWR VGND _03680_ sg13g2_nand3_1
X_09948_ _03651_ _03650_ VPWR VGND _03681_ sg13g2_nand2b_1
X_09949_ _03649_ _03678_ _03681_ VPWR VGND _03682_ sg13g2_nand3b_1
X_09950_ _01599_ _03636_ VPWR VGND _03683_ sg13g2_xor2_1
X_09951_ _01713_ _03636_ VPWR VGND _03684_ sg13g2_nand2_1
X_09952_ _02029_ _03667_ _03684_ VPWR VGND _03685_ sg13g2_a21oi_1
X_09953_ _03667_ _03683_ _03685_ VPWR VGND _03686_ sg13g2_a21oi_1
X_09954_ _03609_ _01907_ VPWR VGND _03687_ sg13g2_xor2_1
X_09955_ _03612_ _03635_ VPWR VGND _03688_ sg13g2_xnor2_1
X_09956_ _01858_ _03688_ VPWR VGND _03689_ sg13g2_xor2_1
X_09957_ _03628_ _03629_ VPWR VGND _03690_ sg13g2_nand2_1
X_09958_ _01667_ _03630_ VPWR VGND _03691_ sg13g2_xnor2_1
X_09959_ _03690_ _03691_ VPWR VGND _03692_ sg13g2_xnor2_1
X_09960_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[24]\ VPWR VGND _03693_ sg13g2_inv_1
X_09961_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[22]\ VPWR VGND _03694_ sg13g2_inv_1
X_09962_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ VPWR VGND _03695_ sg13g2_inv_1
X_09963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[20]\ VPWR VGND _03696_ sg13g2_inv_1
X_09964_ _01791_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ VPWR VGND _03697_ sg13g2_nand2b_1
X_09965_ _03696_ _03697_ VPWR VGND _03698_ sg13g2_nand2_1
X_09966_ _03696_ _03697_ VPWR VGND _03699_ sg13g2_nor2_1
X_09967_ _01965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ _03698_ _01796_ _03699_ VPWR 
+ VGND
+ _03700_ sg13g2_a221oi_1
X_09968_ _01801_ _03694_ _03695_ _01787_ _03700_ VPWR 
+ VGND
+ _03701_ sg13g2_a221oi_1
X_09969_ _01963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ VPWR VGND _03702_ sg13g2_nand2_1
X_09970_ _01801_ _03694_ _03702_ VPWR VGND _03703_ sg13g2_o21ai_1
X_09971_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ _01783_ VPWR VGND _03704_ sg13g2_nand2b_1
X_09972_ _03701_ _03703_ _03704_ VPWR VGND _03705_ sg13g2_o21ai_1
X_09973_ _03693_ _03705_ _01809_ VPWR VGND _03706_ sg13g2_o21ai_1
X_09974_ _03693_ _03705_ VPWR VGND _03707_ sg13g2_nand2_1
X_09975_ _01767_ _03617_ VPWR VGND _03708_ sg13g2_xnor2_1
X_09976_ _03132_ _03708_ VPWR VGND _03709_ sg13g2_xor2_1
X_09977_ _03616_ _01774_ VPWR VGND _03710_ sg13g2_xor2_1
X_09978_ _03706_ _03707_ _03709_ _01956_ _03710_ VPWR 
+ VGND
+ _03711_ sg13g2_a221oi_1
X_09979_ _03616_ _03109_ VPWR VGND _03712_ sg13g2_nand2b_1
X_09980_ _01819_ _03616_ _03107_ VPWR VGND _03713_ sg13g2_nand3_1
X_09981_ _01832_ VPWR VGND _03714_ sg13g2_inv_1
X_09982_ _01834_ _03616_ _01761_ VPWR VGND _03715_ sg13g2_o21ai_1
X_09983_ _01834_ _03616_ _01761_ VPWR VGND _03716_ sg13g2_a21oi_1
X_09984_ _03714_ _03715_ _03716_ VPWR VGND _03717_ sg13g2_a21oi_1
X_09985_ _03713_ _03717_ _03708_ VPWR VGND _03718_ sg13g2_mux2_1
X_09986_ _03613_ _01750_ VPWR VGND _03719_ sg13g2_xnor2_1
X_09987_ _03719_ VPWR VGND _03720_ sg13g2_inv_1
X_09988_ _01735_ _03624_ _03720_ VPWR VGND _03721_ sg13g2_nor3_1
X_09989_ _03625_ _01735_ _03624_ VPWR VGND _03722_ sg13g2_nand3b_1
X_09990_ _01744_ _03625_ VPWR VGND _03723_ sg13g2_nand2_1
X_09991_ _03722_ _03723_ _03719_ VPWR VGND _03724_ sg13g2_a21oi_1
X_09992_ _03721_ _03724_ _02687_ VPWR VGND _03725_ sg13g2_o21ai_1
X_09993_ _01758_ _03618_ _03619_ VPWR VGND _03726_ sg13g2_a21oi_1
X_09994_ _01753_ _03614_ VPWR VGND _03727_ sg13g2_xnor2_1
X_09995_ _03726_ _03727_ VPWR VGND _03728_ sg13g2_xnor2_1
X_09996_ _01814_ _03728_ VPWR VGND _03729_ sg13g2_nand2_1
X_09997_ _03712_ _03718_ _03725_ _03729_ VPWR VGND 
+ _03730_
+ sg13g2_nand4_1
X_09998_ _01738_ _03625_ _03624_ VPWR VGND _03731_ sg13g2_o21ai_1
X_09999_ _01738_ _03624_ VPWR VGND _03732_ sg13g2_nor2_1
X_10000_ _01744_ _03731_ _03732_ VPWR VGND _03733_ sg13g2_a21oi_1
X_10001_ _01989_ _03728_ VPWR VGND _03734_ sg13g2_xnor2_1
X_10002_ _03734_ _03729_ VPWR VGND _03735_ sg13g2_and2_1
X_10003_ _01744_ _03622_ VPWR VGND _03736_ sg13g2_nor2_1
X_10004_ _03615_ _03621_ VPWR VGND _03737_ sg13g2_nor2_1
X_10005_ _01738_ _03737_ VPWR VGND _03738_ sg13g2_nand2_1
X_10006_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[9]\ VPWR VGND _03739_ sg13g2_xor2_1
X_10007_ _03736_ _03738_ _03739_ _03737_ _03719_ VPWR 
+ VGND
+ _03740_ sg13g2_a221oi_1
X_10008_ _03719_ _03733_ _03725_ _03735_ _03740_ VPWR 
+ VGND
+ _03741_ sg13g2_a221oi_1
X_10009_ _03711_ _03730_ _03741_ VPWR VGND _03742_ sg13g2_o21ai_1
X_10010_ _01729_ _03613_ VPWR VGND _03743_ sg13g2_xor2_1
X_10011_ _03627_ _03743_ VPWR VGND _03744_ sg13g2_xnor2_1
X_10012_ _01727_ _03744_ VPWR VGND _03745_ sg13g2_nand2_1
X_10013_ _03692_ _03742_ _03745_ VPWR VGND _03746_ sg13g2_nand3_1
X_10014_ _01850_ _03742_ _03745_ VPWR VGND _03747_ sg13g2_nand3_1
X_10015_ _02731_ _03692_ VPWR VGND _03748_ sg13g2_nand2_1
X_10016_ _03689_ _03746_ _03747_ _03748_ VPWR VGND 
+ _03749_
+ sg13g2_nand4_1
X_10017_ _01725_ _03665_ _03683_ VPWR VGND _03750_ sg13g2_nand3_1
X_10018_ _02572_ _03688_ _03750_ VPWR VGND _03751_ sg13g2_o21ai_1
X_10019_ _01951_ _02572_ VPWR VGND _03752_ sg13g2_nor2_1
X_10020_ _03611_ _03683_ VPWR VGND _03753_ sg13g2_nor2_1
X_10021_ _03611_ _03683_ VPWR VGND _03754_ sg13g2_nand2_1
X_10022_ _03632_ _03633_ _03754_ VPWR VGND _03755_ sg13g2_a21oi_1
X_10023_ _03635_ _03753_ _03755_ VPWR VGND _03756_ sg13g2_a21oi_1
X_10024_ _03663_ _03683_ VPWR VGND _03757_ sg13g2_or2_1
X_10025_ _03756_ _03757_ _02029_ VPWR VGND _03758_ sg13g2_a21oi_1
X_10026_ _01951_ _03751_ _03752_ _03688_ _03758_ VPWR 
+ VGND
+ _03759_ sg13g2_a221oi_1
X_10027_ _01946_ _02029_ _03663_ _03665_ _03636_ VPWR 
+ VGND
+ _03760_ sg13g2_a221oi_1
X_10028_ _03636_ _03667_ _02032_ VPWR VGND _03761_ sg13g2_a21oi_1
X_10029_ _03687_ _03760_ _03761_ VPWR VGND _03762_ sg13g2_nor3_1
X_10030_ _03686_ _03687_ _03749_ _03759_ _03762_ VPWR 
+ VGND
+ _03763_ sg13g2_a221oi_1
X_10031_ _03680_ _03682_ _03763_ VPWR VGND _03764_ sg13g2_a21oi_1
X_10032_ _02036_ _03678_ VPWR VGND _03765_ sg13g2_nand2_1
X_10033_ _02036_ _03681_ VPWR VGND _03766_ sg13g2_nand2_1
X_10034_ _02036_ _03679_ VPWR VGND _03767_ sg13g2_nand2_1
X_10035_ _03766_ _03767_ _03649_ VPWR VGND _03768_ sg13g2_mux2_1
X_10036_ _01880_ _03768_ VPWR VGND _03769_ sg13g2_and2_1
X_10037_ _03763_ _03765_ _03769_ VPWR VGND _03770_ sg13g2_o21ai_1
X_10038_ _03764_ _03770_ _03396_ VPWR VGND _03771_ sg13g2_o21ai_1
X_10039_ _02064_ _03607_ VPWR VGND _03772_ sg13g2_xnor2_1
X_10040_ _03652_ _03772_ VPWR VGND _03773_ sg13g2_xnor2_1
X_10041_ _03763_ _03765_ VPWR VGND _03774_ sg13g2_nor2_1
X_10042_ _01880_ _03768_ VPWR VGND _03775_ sg13g2_nand2b_1
X_10043_ _03774_ _03764_ _03773_ _03775_ VPWR VGND 
+ _03776_
+ sg13g2_nor4_1
X_10044_ _03771_ _03773_ _03776_ VPWR VGND _03777_ sg13g2_a21o_1
X_10045_ _01897_ _03659_ _03661_ _03777_ VPWR VGND 
+ _03778_
+ sg13g2_nand4_1
X_10046_ _01897_ _03661_ VPWR VGND _03779_ sg13g2_nor2_1
X_10047_ _03659_ _03777_ _03779_ VPWR VGND _03780_ sg13g2_nand3_1
X_10048_ _02086_ _03659_ _03661_ VPWR VGND _03781_ sg13g2_nand3_1
X_10049_ _02108_ _03778_ _03780_ _03781_ VPWR VGND 
+ _03782_
+ sg13g2_nand4_1
X_10050_ _01901_ _02448_ VPWR VGND _03783_ sg13g2_nand2_1
X_10051_ _03606_ _03782_ _03783_ VPWR VGND _00453_ sg13g2_o21ai_1
X_10052_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2073_o[1]\ VPWR VGND _03784_ sg13g2_buf_1
X_10053_ _03784_ VPWR VGND _03785_ sg13g2_inv_1
X_10054_ _02771_ _02448_ VPWR VGND _03786_ sg13g2_nand2_1
X_10055_ _03785_ _03782_ _03786_ VPWR VGND _00454_ sg13g2_o21ai_1
X_10056_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2076_o[0]\ VPWR VGND _03787_ sg13g2_buf_1
X_10057_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[17]\ VPWR VGND _03788_ sg13g2_buf_1
X_10058_ _03788_ VPWR VGND _03789_ sg13g2_inv_1
X_10059_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2078_o\ VPWR VGND _03790_ sg13g2_inv_1
X_10060_ _03789_ _03790_ VPWR VGND _03791_ sg13g2_nor2_1
X_10061_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[13]\ VPWR VGND _03792_ sg13g2_buf_1
X_10062_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[11]\ VPWR VGND _03793_ sg13g2_inv_1
X_10063_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[10]\ VPWR VGND _03794_ sg13g2_buf_1
X_10064_ _03794_ VPWR VGND _03795_ sg13g2_inv_1
X_10065_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[9]\ VPWR VGND _03796_ sg13g2_buf_1
X_10066_ _03796_ VPWR VGND _03797_ sg13g2_inv_1
X_10067_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[8]\ VPWR VGND _03798_ sg13g2_buf_1
X_10068_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[6]\ VPWR VGND _03799_ sg13g2_buf_1
X_10069_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[7]\ VPWR VGND _03800_ sg13g2_buf_1
X_10070_ _01609_ _03799_ _03800_ VPWR VGND _03801_ sg13g2_a21o_1
X_10071_ _01609_ _03800_ _03799_ VPWR VGND _03802_ sg13g2_and3_1
X_10072_ _01614_ _03801_ _03802_ VPWR VGND _03803_ sg13g2_a21o_1
X_10073_ _03803_ VPWR VGND _03804_ sg13g2_buf_1
X_10074_ _03798_ _03804_ VPWR VGND _03805_ sg13g2_nand2_1
X_10075_ _03798_ _03804_ _01753_ VPWR VGND _03806_ sg13g2_o21ai_1
X_10076_ _03797_ _03805_ _03806_ VPWR VGND _03807_ sg13g2_nand3_1
X_10077_ _03807_ VPWR VGND _03808_ sg13g2_buf_1
X_10078_ _03805_ _03806_ _03797_ VPWR VGND _03809_ sg13g2_a21oi_1
X_10079_ _01735_ _03808_ _03809_ VPWR VGND _03810_ sg13g2_a21oi_1
X_10080_ _03795_ _03810_ VPWR VGND _03811_ sg13g2_nor2_1
X_10081_ _03795_ _03810_ _01628_ VPWR VGND _03812_ sg13g2_a21oi_1
X_10082_ _03811_ _03812_ _01666_ VPWR VGND _03813_ sg13g2_o21ai_1
X_10083_ _01666_ _03811_ _03812_ VPWR VGND _03814_ sg13g2_nor3_1
X_10084_ _03793_ _03813_ _03814_ VPWR VGND _03815_ sg13g2_a21oi_1
X_10085_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[12]\ VPWR VGND _03816_ sg13g2_buf_1
X_10086_ _03816_ VPWR VGND _03817_ sg13g2_inv_1
X_10087_ _02419_ _03817_ VPWR VGND _03818_ sg13g2_nand2_1
X_10088_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[14]\ VPWR VGND _03819_ sg13g2_buf_1
X_10089_ _01672_ _03819_ VPWR VGND _03820_ sg13g2_nand2_1
X_10090_ _02419_ _03817_ _03820_ VPWR VGND _03821_ sg13g2_o21ai_1
X_10091_ _01713_ _03792_ _03815_ _03818_ _03821_ VPWR 
+ VGND
+ _03822_ sg13g2_a221oi_1
X_10092_ _01712_ _03792_ VPWR VGND _03823_ sg13g2_nor2_1
X_10093_ _03823_ _03820_ VPWR VGND _03824_ sg13g2_nand2_1
X_10094_ _01706_ _03819_ _03824_ VPWR VGND _03825_ sg13g2_o21ai_1
X_10095_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[15]\ VPWR VGND _03826_ sg13g2_inv_1
X_10096_ _03822_ _03825_ _03826_ VPWR VGND _03827_ sg13g2_o21ai_1
X_10097_ _03826_ _03822_ _03825_ VPWR VGND _03828_ sg13g2_nor3_1
X_10098_ _01877_ _03827_ _03828_ VPWR VGND _03829_ sg13g2_a21oi_1
X_10099_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[16]\ VPWR VGND _03830_ sg13g2_buf_1
X_10100_ _01682_ _03830_ VPWR VGND _03831_ sg13g2_nand2_1
X_10101_ _01682_ _03830_ VPWR VGND _03832_ sg13g2_nor2_1
X_10102_ _03829_ _03831_ _03832_ VPWR VGND _03833_ sg13g2_a21oi_1
X_10103_ _03789_ _03791_ _03833_ VPWR VGND _03834_ sg13g2_mux2_1
X_10104_ _03789_ _03833_ VPWR VGND _03835_ sg13g2_xnor2_1
X_10105_ _03790_ _02289_ _02290_ VPWR VGND _03836_ sg13g2_o21ai_1
X_10106_ _02292_ _03834_ _03835_ _03836_ VPWR VGND 
+ _03837_
+ sg13g2_a22oi_1
X_10107_ _02419_ _03817_ VPWR VGND _03838_ sg13g2_nor2_1
X_10108_ _02419_ _03817_ _03793_ _03813_ _03814_ VPWR 
+ VGND
+ _03839_ sg13g2_a221oi_1
X_10109_ _03792_ _03838_ _03839_ VPWR VGND _03840_ sg13g2_or3_1
X_10110_ _03819_ _01908_ VPWR VGND _03841_ sg13g2_xnor2_1
X_10111_ _03840_ _03841_ _01912_ VPWR VGND _03842_ sg13g2_nand3b_1
X_10112_ _03838_ _03839_ _03792_ VPWR VGND _03843_ sg13g2_o21ai_1
X_10113_ _03819_ _01907_ VPWR VGND _03844_ sg13g2_xor2_1
X_10114_ _01947_ _03840_ _03843_ _03844_ VPWR VGND 
+ _03845_
+ sg13g2_nand4_1
X_10115_ _03843_ _03844_ _01912_ VPWR VGND _03846_ sg13g2_nand3b_1
X_10116_ _03842_ _03845_ _03846_ VPWR VGND _03847_ sg13g2_nand3_1
X_10117_ _03838_ _03818_ VPWR VGND _03848_ sg13g2_nor2b_1
X_10118_ _03815_ _03848_ VPWR VGND _03849_ sg13g2_xnor2_1
X_10119_ _01735_ _03808_ _03809_ VPWR VGND _03850_ sg13g2_a21o_1
X_10120_ _03850_ VPWR VGND _03851_ sg13g2_buf_1
X_10121_ _03794_ _03851_ VPWR VGND _03852_ sg13g2_nand2_1
X_10122_ _03794_ _03851_ _01729_ VPWR VGND _03853_ sg13g2_o21ai_1
X_10123_ _03852_ _03853_ _03793_ VPWR VGND _03854_ sg13g2_a21oi_1
X_10124_ _03793_ _03852_ _03853_ VPWR VGND _03855_ sg13g2_nand3_1
X_10125_ _01850_ _03854_ _03855_ VPWR VGND _03856_ sg13g2_o21ai_1
X_10126_ _01850_ _03855_ VPWR VGND _03857_ sg13g2_nor2_1
X_10127_ _02018_ _03856_ _03857_ VPWR VGND _03858_ sg13g2_a21oi_1
X_10128_ _03816_ _01858_ VPWR VGND _03859_ sg13g2_xnor2_1
X_10129_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[43]\ VPWR VGND _03860_ sg13g2_inv_1
X_10130_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[42]\ VPWR VGND _03861_ sg13g2_inv_1
X_10131_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[40]\ VPWR VGND _03862_ sg13g2_inv_1
X_10132_ _01788_ _03862_ VPWR VGND _03863_ sg13g2_nor2_1
X_10133_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ VPWR VGND _03864_ sg13g2_nor2b_1
X_10134_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _03864_ VPWR VGND _03865_ sg13g2_nand2_1
X_10135_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _03864_ _01796_ VPWR VGND _03866_ sg13g2_o21ai_1
X_10136_ _01788_ _03862_ _03865_ _03866_ VPWR VGND 
+ _03867_
+ sg13g2_a22oi_1
X_10137_ _03863_ _03867_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ VPWR VGND _03868_ sg13g2_o21ai_1
X_10138_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _03863_ _03867_ VPWR VGND _03869_ sg13g2_nor3_1
X_10139_ _01783_ _03861_ _03868_ _01803_ _03869_ VPWR 
+ VGND
+ _03870_ sg13g2_a221oi_1
X_10140_ _01964_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[42]\ _03870_ VPWR VGND _03871_ sg13g2_a21oi_1
X_10141_ _03860_ _03871_ _01810_ VPWR VGND _03872_ sg13g2_o21ai_1
X_10142_ _03860_ _03871_ VPWR VGND _03873_ sg13g2_nand2_1
X_10143_ _03798_ _01756_ VPWR VGND _03874_ sg13g2_xnor2_1
X_10144_ _01761_ _03802_ _03801_ VPWR VGND _03875_ sg13g2_o21ai_1
X_10145_ _01780_ _03875_ VPWR VGND _03876_ sg13g2_nand2_1
X_10146_ _01841_ _03801_ _03876_ VPWR VGND _03877_ sg13g2_o21ai_1
X_10147_ _01832_ _01840_ _03799_ VPWR VGND _03878_ sg13g2_nand3_1
X_10148_ _01759_ _03800_ _03878_ VPWR VGND _03879_ sg13g2_nand3_1
X_10149_ _01818_ _03799_ VPWR VGND _03880_ sg13g2_nand2_1
X_10150_ _01767_ _03800_ VPWR VGND _03881_ sg13g2_xor2_1
X_10151_ _03880_ _03881_ VPWR VGND _03882_ sg13g2_nand2b_1
X_10152_ _03879_ _03882_ _03874_ VPWR VGND _03883_ sg13g2_a21oi_1
X_10153_ _03874_ _03877_ _03883_ VPWR VGND _03884_ sg13g2_a21o_1
X_10154_ _03799_ _01774_ VPWR VGND _03885_ sg13g2_xnor2_1
X_10155_ _03884_ _03885_ VPWR VGND _03886_ sg13g2_nand2_1
X_10156_ _03872_ _03873_ _03886_ VPWR VGND _03887_ sg13g2_a21oi_1
X_10157_ _03805_ _03806_ VPWR VGND _03888_ sg13g2_nand2_1
X_10158_ _01740_ _03796_ VPWR VGND _03889_ sg13g2_xor2_1
X_10159_ _03888_ _03889_ VPWR VGND _03890_ sg13g2_xor2_1
X_10160_ _03880_ _03881_ VPWR VGND _03891_ sg13g2_xnor2_1
X_10161_ _01819_ _03799_ VPWR VGND _03892_ sg13g2_or2_1
X_10162_ _03880_ _03892_ _01983_ VPWR VGND _03893_ sg13g2_a21o_1
X_10163_ _01956_ _03891_ _03893_ VPWR VGND _03894_ sg13g2_o21ai_1
X_10164_ _01990_ _03798_ VPWR VGND _03895_ sg13g2_xor2_1
X_10165_ _03804_ _03895_ VPWR VGND _03896_ sg13g2_xnor2_1
X_10166_ _03884_ _03894_ _03896_ _01998_ VPWR VGND 
+ _03897_
+ sg13g2_a22oi_1
X_10167_ _01812_ _03890_ _03897_ VPWR VGND _03898_ sg13g2_o21ai_1
X_10168_ _01740_ _03796_ VPWR VGND _03899_ sg13g2_nand2_1
X_10169_ _01739_ _03888_ _03899_ VPWR VGND _03900_ sg13g2_a21oi_1
X_10170_ _03888_ _03889_ _03900_ VPWR VGND _03901_ sg13g2_a21oi_1
X_10171_ _03794_ _01750_ VPWR VGND _03902_ sg13g2_xnor2_1
X_10172_ _01738_ _03809_ _03808_ VPWR VGND _03903_ sg13g2_o21ai_1
X_10173_ _01744_ _03903_ VPWR VGND _03904_ sg13g2_and2_1
X_10174_ _01812_ _03808_ VPWR VGND _03905_ sg13g2_nor2_1
X_10175_ _03904_ _03905_ _03902_ VPWR VGND _03906_ sg13g2_o21ai_1
X_10176_ _03901_ _03902_ _03906_ VPWR VGND _03907_ sg13g2_o21ai_1
X_10177_ _03887_ _03898_ _03907_ VPWR VGND _03908_ sg13g2_o21ai_1
X_10178_ _01730_ _03794_ VPWR VGND _03909_ sg13g2_xor2_1
X_10179_ _03851_ _03909_ VPWR VGND _03910_ sg13g2_xnor2_1
X_10180_ _03852_ _03853_ VPWR VGND _03911_ sg13g2_nand2_1
X_10181_ _01667_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[11]\ VPWR VGND _03912_ sg13g2_xor2_1
X_10182_ _03911_ _03912_ VPWR VGND _03913_ sg13g2_xnor2_1
X_10183_ _02250_ _03910_ _03913_ _02014_ VPWR VGND 
+ _03914_
+ sg13g2_a22oi_1
X_10184_ _02018_ _03793_ VPWR VGND _03915_ sg13g2_nor2_1
X_10185_ _01850_ _03911_ VPWR VGND _03916_ sg13g2_nand2_1
X_10186_ _03915_ _03916_ _03912_ _03911_ _03859_ VPWR 
+ VGND
+ _03917_ sg13g2_a221oi_1
X_10187_ _03858_ _03859_ _03908_ _03914_ _03917_ VPWR 
+ VGND
+ _03918_ sg13g2_a221oi_1
X_10188_ _01722_ _03849_ _03918_ VPWR VGND _03919_ sg13g2_a21o_1
X_10189_ _01947_ _03792_ _03844_ VPWR VGND _03920_ sg13g2_nand3_1
X_10190_ _01946_ _03792_ _03816_ _01951_ _03839_ VPWR 
+ VGND
+ _03921_ sg13g2_a221oi_1
X_10191_ _03823_ _03921_ _03841_ VPWR VGND _03922_ sg13g2_o21ai_1
X_10192_ _03920_ _03922_ _02029_ VPWR VGND _03923_ sg13g2_a21oi_1
X_10193_ _01913_ _03847_ _03919_ _03923_ VPWR VGND 
+ _03924_
+ sg13g2_a22oi_1
X_10194_ _03823_ _03921_ VPWR VGND _03925_ sg13g2_nor2_1
X_10195_ _01872_ _03819_ VPWR VGND _03926_ sg13g2_xor2_1
X_10196_ _03925_ _03926_ VPWR VGND _03927_ sg13g2_xnor2_1
X_10197_ _03847_ _03919_ _03927_ _02048_ VPWR VGND 
+ _03928_
+ sg13g2_a22oi_1
X_10198_ _03924_ _03928_ VPWR VGND _03929_ sg13g2_nand2_1
X_10199_ _02343_ _03830_ VPWR VGND _03930_ sg13g2_xnor2_1
X_10200_ _03829_ _03930_ VPWR VGND _03931_ sg13g2_xnor2_1
X_10201_ _03847_ _03919_ _03927_ _02048_ _01887_ VPWR 
+ VGND
+ _03932_ sg13g2_a221oi_1
X_10202_ _03822_ _03825_ VPWR VGND _03933_ sg13g2_nor2_1
X_10203_ _02044_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[15]\ VPWR VGND _03934_ sg13g2_xnor2_1
X_10204_ _03933_ _03934_ VPWR VGND _03935_ sg13g2_xnor2_1
X_10205_ _03924_ _03932_ _03935_ VPWR VGND _03936_ sg13g2_a21oi_1
X_10206_ _01887_ _03929_ _03931_ _01890_ _03936_ VPWR 
+ VGND
+ _03937_ sg13g2_a221oi_1
X_10207_ _02278_ _02752_ _03931_ VPWR VGND _03938_ sg13g2_mux2_1
X_10208_ _03837_ _03937_ _03938_ VPWR VGND _03939_ sg13g2_nor3_1
X_10209_ _02089_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2078_o\ _03835_ VPWR VGND _03940_ sg13g2_nand3_1
X_10210_ _02088_ _03788_ _03833_ VPWR VGND _03941_ sg13g2_nor3_1
X_10211_ _01697_ _03788_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2078_o\ _03833_ VPWR VGND 
+ _03942_
+ sg13g2_nand4_1
X_10212_ _03941_ _03942_ VPWR VGND _03943_ sg13g2_nor2b_1
X_10213_ _03940_ _03943_ _01895_ VPWR VGND _03944_ sg13g2_a21oi_1
X_10214_ _02589_ _03939_ _03944_ VPWR VGND _03945_ sg13g2_nor3_1
X_10215_ _03606_ _01903_ VPWR VGND _03946_ sg13g2_nor2_1
X_10216_ _03787_ _03945_ _03946_ VPWR VGND _00455_ sg13g2_a21o_1
X_10217_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2076_o[1]\ VPWR VGND _03947_ sg13g2_buf_1
X_10218_ _03785_ _01903_ VPWR VGND _03948_ sg13g2_nor2_1
X_10219_ _03947_ _03945_ _03948_ VPWR VGND _00456_ sg13g2_a21o_1
X_10220_ _03787_ _02924_ VPWR VGND _03949_ sg13g2_nand2_1
X_10221_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2079_o[0]\ VPWR VGND _03950_ sg13g2_buf_1
X_10222_ _03950_ _01903_ VPWR VGND _03951_ sg13g2_nand2_1
X_10223_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[12]\ VPWR VGND _03952_ sg13g2_buf_1
X_10224_ _03952_ VPWR VGND _03953_ sg13g2_inv_1
X_10225_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[11]\ VPWR VGND _03954_ sg13g2_inv_1
X_10226_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[10]\ VPWR VGND _03955_ sg13g2_buf_1
X_10227_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[8]\ VPWR VGND _03956_ sg13g2_buf_1
X_10228_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[6]\ VPWR VGND _03957_ sg13g2_buf_1
X_10229_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[7]\ VPWR VGND _03958_ sg13g2_buf_1
X_10230_ _01763_ _03957_ _03958_ VPWR VGND _03959_ sg13g2_a21o_1
X_10231_ _03959_ VPWR VGND _03960_ sg13g2_buf_1
X_10232_ _01763_ _03958_ _03957_ VPWR VGND _03961_ sg13g2_and3_1
X_10233_ _03961_ VPWR VGND _03962_ sg13g2_buf_1
X_10234_ _01619_ _03956_ _03960_ _01758_ _03962_ VPWR 
+ VGND
+ _03963_ sg13g2_a221oi_1
X_10235_ _01753_ _03956_ VPWR VGND _03964_ sg13g2_nor2_1
X_10236_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[9]\ VPWR VGND _03965_ sg13g2_inv_1
X_10237_ _03963_ _03964_ _03965_ VPWR VGND _03966_ sg13g2_o21ai_1
X_10238_ _03965_ _03963_ _03964_ VPWR VGND _03967_ sg13g2_nor3_1
X_10239_ _01735_ _03966_ _03967_ VPWR VGND _03968_ sg13g2_a21o_1
X_10240_ _03968_ VPWR VGND _03969_ sg13g2_buf_1
X_10241_ _03955_ _03969_ VPWR VGND _03970_ sg13g2_nand2_1
X_10242_ _03955_ _03969_ _01729_ VPWR VGND _03971_ sg13g2_o21ai_1
X_10243_ _03954_ _03970_ _03971_ VPWR VGND _03972_ sg13g2_nand3_1
X_10244_ _03970_ _03971_ _03954_ VPWR VGND _03973_ sg13g2_a21oi_1
X_10245_ _01853_ _03972_ _03973_ VPWR VGND _03974_ sg13g2_a21oi_1
X_10246_ _03974_ VPWR VGND _03975_ sg13g2_inv_1
X_10247_ _03952_ _03975_ _01951_ VPWR VGND _03976_ sg13g2_a21oi_1
X_10248_ _03953_ _03974_ _03976_ VPWR VGND _03977_ sg13g2_a21oi_1
X_10249_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[13]\ VPWR VGND _03978_ sg13g2_buf_1
X_10250_ _01947_ _03978_ VPWR VGND _03979_ sg13g2_xnor2_1
X_10251_ _03977_ _03979_ VPWR VGND _03980_ sg13g2_xnor2_1
X_10252_ _01729_ _03955_ VPWR VGND _03981_ sg13g2_xor2_1
X_10253_ _03969_ _03981_ VPWR VGND _03982_ sg13g2_xnor2_1
X_10254_ _03982_ VPWR VGND _03983_ sg13g2_buf_1
X_10255_ _03963_ _03964_ VPWR VGND _03984_ sg13g2_nor2_1
X_10256_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[9]\ VPWR VGND _03985_ sg13g2_xnor2_1
X_10257_ _03984_ _03985_ VPWR VGND _03986_ sg13g2_xnor2_1
X_10258_ _01748_ _03983_ _03986_ VPWR VGND _03987_ sg13g2_or3_1
X_10259_ _01748_ _01812_ _03983_ VPWR VGND _03988_ sg13g2_or3_1
X_10260_ _01959_ _03960_ _03962_ VPWR VGND _03989_ sg13g2_a21oi_1
X_10261_ _01990_ _03956_ VPWR VGND _03990_ sg13g2_xnor2_1
X_10262_ _03989_ _03990_ VPWR VGND _03991_ sg13g2_xnor2_1
X_10263_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[62]\ VPWR VGND _03992_ sg13g2_inv_1
X_10264_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[60]\ VPWR VGND _03993_ sg13g2_inv_1
X_10265_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[59]\ VPWR VGND _03994_ sg13g2_inv_1
X_10266_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[58]\ VPWR VGND _03995_ sg13g2_inv_1
X_10267_ _01970_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ VPWR VGND _03996_ sg13g2_nand2b_1
X_10268_ _03995_ _03996_ VPWR VGND _03997_ sg13g2_nand2_1
X_10269_ _03995_ _03996_ VPWR VGND _03998_ sg13g2_nor2_1
X_10270_ _01966_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[59]\ _03997_ _01797_ _03998_ VPWR 
+ VGND
+ _03999_ sg13g2_a221oi_1
X_10271_ _01802_ _03993_ _03994_ _02382_ _03999_ VPWR 
+ VGND
+ _04000_ sg13g2_a221oi_1
X_10272_ _01964_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ VPWR VGND _04001_ sg13g2_nand2_1
X_10273_ _01802_ _03993_ _04001_ VPWR VGND _04002_ sg13g2_o21ai_1
X_10274_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ _01783_ VPWR VGND _04003_ sg13g2_nand2b_1
X_10275_ _04000_ _04002_ _04003_ VPWR VGND _04004_ sg13g2_o21ai_1
X_10276_ _01810_ _03992_ _04004_ VPWR VGND _04005_ sg13g2_a21o_1
X_10277_ _01818_ _03957_ VPWR VGND _04006_ sg13g2_nand2_1
X_10278_ _01758_ _03958_ VPWR VGND _04007_ sg13g2_xnor2_1
X_10279_ _01818_ _01760_ _03957_ VPWR VGND _04008_ sg13g2_nand3_1
X_10280_ _01767_ _03958_ _04008_ VPWR VGND _04009_ sg13g2_nand3_1
X_10281_ _04006_ _04007_ _04009_ VPWR VGND _04010_ sg13g2_o21ai_1
X_10282_ _03956_ _01756_ VPWR VGND _04011_ sg13g2_xnor2_1
X_10283_ _01760_ _03962_ _03960_ VPWR VGND _04012_ sg13g2_o21ai_1
X_10284_ _01761_ _03960_ VPWR VGND _04013_ sg13g2_nor2_1
X_10285_ _01780_ _04012_ _04013_ VPWR VGND _04014_ sg13g2_a21oi_1
X_10286_ _04011_ _04014_ VPWR VGND _04015_ sg13g2_nand2_1
X_10287_ _04010_ _04011_ _04015_ VPWR VGND _04016_ sg13g2_o21ai_1
X_10288_ _03957_ _01774_ VPWR VGND _04017_ sg13g2_xnor2_1
X_10289_ _01810_ _03992_ _04017_ VPWR VGND _04018_ sg13g2_o21ai_1
X_10290_ _04016_ _04018_ VPWR VGND _04019_ sg13g2_nor2_1
X_10291_ _01957_ _03957_ VPWR VGND _04020_ sg13g2_xnor2_1
X_10292_ _04006_ _04007_ VPWR VGND _04021_ sg13g2_xnor2_1
X_10293_ _01827_ _04020_ _04021_ _02548_ VPWR VGND 
+ _04022_
+ sg13g2_a22oi_1
X_10294_ _04016_ _04022_ VPWR VGND _04023_ sg13g2_nor2_1
X_10295_ _01998_ _03991_ _04005_ _04019_ _04023_ VPWR 
+ VGND
+ _04024_ sg13g2_a221oi_1
X_10296_ _03987_ _03988_ _04024_ VPWR VGND _04025_ sg13g2_a21o_1
X_10297_ _03986_ VPWR VGND _04026_ sg13g2_inv_1
X_10298_ _01748_ _03983_ _04026_ VPWR VGND _04027_ sg13g2_nand3_1
X_10299_ _02254_ _01739_ VPWR VGND _04028_ sg13g2_nor2_1
X_10300_ _04028_ _03983_ VPWR VGND _04029_ sg13g2_nand2_1
X_10301_ _04027_ _04029_ _04024_ VPWR VGND _04030_ sg13g2_a21o_1
X_10302_ _01748_ _01812_ _03983_ _03986_ VPWR VGND 
+ _04031_
+ sg13g2_nor4_1
X_10303_ _04028_ _03983_ _04026_ VPWR VGND _04032_ sg13g2_nand3_1
X_10304_ _04031_ _04032_ VPWR VGND _04033_ sg13g2_nand2b_1
X_10305_ _01727_ _03983_ _04033_ VPWR VGND _04034_ sg13g2_a21oi_1
X_10306_ _04025_ _04030_ _04034_ VPWR VGND _04035_ sg13g2_nand3_1
X_10307_ _03970_ _03971_ VPWR VGND _04036_ sg13g2_nand2_1
X_10308_ _01853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[11]\ VPWR VGND _04037_ sg13g2_xor2_1
X_10309_ _04036_ _04037_ VPWR VGND _04038_ sg13g2_xnor2_1
X_10310_ _02015_ _04035_ _04038_ VPWR VGND _04039_ sg13g2_a21oi_1
X_10311_ _02731_ _04025_ _04030_ _04034_ VPWR VGND 
+ _04040_
+ sg13g2_nand4_1
X_10312_ _01856_ _04040_ VPWR VGND _04041_ sg13g2_nand2_1
X_10313_ _04039_ _04041_ _02572_ VPWR VGND _04042_ sg13g2_o21ai_1
X_10314_ _01951_ _03952_ VPWR VGND _04043_ sg13g2_xor2_1
X_10315_ _03974_ _04043_ VPWR VGND _04044_ sg13g2_xnor2_1
X_10316_ _02571_ _04040_ VPWR VGND _04045_ sg13g2_nand2_1
X_10317_ _04039_ _04045_ _04044_ VPWR VGND _04046_ sg13g2_o21ai_1
X_10318_ _04042_ _04044_ _04046_ VPWR VGND _04047_ sg13g2_o21ai_1
X_10319_ _02575_ _03980_ _04047_ VPWR VGND _04048_ sg13g2_o21ai_1
X_10320_ _01711_ _03978_ VPWR VGND _04049_ sg13g2_nand2_1
X_10321_ _03953_ _04049_ VPWR VGND _04050_ sg13g2_nand2_1
X_10322_ _01915_ _04049_ VPWR VGND _04051_ sg13g2_nand2_1
X_10323_ _01667_ _03972_ _04050_ _04051_ _03973_ VPWR 
+ VGND
+ _04052_ sg13g2_a221oi_1
X_10324_ _01662_ _03952_ VPWR VGND _04053_ sg13g2_nor2_1
X_10325_ _01712_ _03978_ VPWR VGND _04054_ sg13g2_nor2_1
X_10326_ _04049_ _04053_ _04054_ VPWR VGND _04055_ sg13g2_a21oi_1
X_10327_ _04052_ _04055_ VPWR VGND _04056_ sg13g2_nor2b_1
X_10328_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[14]\ VPWR VGND _04057_ sg13g2_buf_1
X_10329_ _04057_ _01908_ VPWR VGND _04058_ sg13g2_xnor2_1
X_10330_ _04057_ VPWR VGND _04059_ sg13g2_inv_1
X_10331_ _04052_ _04055_ VPWR VGND _04060_ sg13g2_nand2b_1
X_10332_ _04060_ VPWR VGND _04061_ sg13g2_buf_2
X_10333_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[15]\ VPWR VGND _04062_ sg13g2_buf_1
X_10334_ _01876_ _04062_ VPWR VGND _04063_ sg13g2_xnor2_1
X_10335_ _02050_ _04063_ VPWR VGND _04064_ sg13g2_xnor2_1
X_10336_ _04059_ _04061_ _04064_ _02037_ VPWR VGND 
+ _04065_
+ sg13g2_a22oi_1
X_10337_ _04057_ _04063_ VPWR VGND _04066_ sg13g2_xnor2_1
X_10338_ _04057_ _04061_ _04066_ _02037_ _01908_ VPWR 
+ VGND
+ _04067_ sg13g2_a221oi_1
X_10339_ _01908_ _04065_ _04067_ VPWR VGND _04068_ sg13g2_a21oi_1
X_10340_ _04056_ _04058_ _03980_ _02575_ _04068_ VPWR 
+ VGND
+ _04069_ sg13g2_a221oi_1
X_10341_ _04048_ _04069_ VPWR VGND _04070_ sg13g2_and2_1
X_10342_ _01658_ _04062_ VPWR VGND _04071_ sg13g2_or2_1
X_10343_ _04071_ VPWR VGND _04072_ sg13g2_buf_1
X_10344_ _04057_ _04056_ _01872_ VPWR VGND _04073_ sg13g2_a21oi_1
X_10345_ _04059_ _04061_ _04073_ VPWR VGND _04074_ sg13g2_a21oi_1
X_10346_ _01595_ _04062_ VPWR VGND _04075_ sg13g2_and2_1
X_10347_ _04075_ VPWR VGND _04076_ sg13g2_buf_1
X_10348_ _04072_ _04074_ _04076_ VPWR VGND _04077_ sg13g2_a21oi_1
X_10349_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[16]\ VPWR VGND _04078_ sg13g2_buf_1
X_10350_ _02343_ _04078_ VPWR VGND _04079_ sg13g2_xor2_1
X_10351_ _04077_ _04079_ VPWR VGND _04080_ sg13g2_xnor2_1
X_10352_ _01873_ _04057_ VPWR VGND _04081_ sg13g2_xor2_1
X_10353_ _04061_ _04081_ _02048_ VPWR VGND _04082_ sg13g2_o21ai_1
X_10354_ _02050_ _04057_ VPWR VGND _04083_ sg13g2_nor2_1
X_10355_ _01703_ _04056_ _02036_ VPWR VGND _04084_ sg13g2_a21oi_1
X_10356_ _02048_ _04061_ VPWR VGND _04085_ sg13g2_nand2_1
X_10357_ _02050_ _04057_ _04085_ VPWR VGND _04086_ sg13g2_nand3_1
X_10358_ _04083_ _04084_ _04086_ VPWR VGND _04087_ sg13g2_o21ai_1
X_10359_ _03229_ _04061_ VPWR VGND _04088_ sg13g2_nand2b_1
X_10360_ _04061_ _04081_ _04083_ _04088_ VPWR VGND 
+ _04089_
+ sg13g2_a22oi_1
X_10361_ _04063_ _04089_ VPWR VGND _04090_ sg13g2_nor2_1
X_10362_ _02037_ _04082_ _04063_ _04087_ _04090_ VPWR 
+ VGND
+ _04091_ sg13g2_a221oi_1
X_10363_ _04091_ VPWR VGND _04092_ sg13g2_inv_1
X_10364_ _03396_ _04080_ _04092_ VPWR VGND _04093_ sg13g2_o21ai_1
X_10365_ _01681_ _04057_ _04072_ VPWR VGND _04094_ sg13g2_nand3_1
X_10366_ _01871_ _01680_ _04072_ VPWR VGND _04095_ sg13g2_nand3_1
X_10367_ _04094_ _04095_ _04061_ VPWR VGND _04096_ sg13g2_a21oi_1
X_10368_ _01681_ _04076_ VPWR VGND _04097_ sg13g2_nand2_1
X_10369_ _04059_ _04095_ _04097_ VPWR VGND _04098_ sg13g2_o21ai_1
X_10370_ _04078_ _04096_ _04098_ VPWR VGND _04099_ sg13g2_nor3_1
X_10371_ _01681_ _04057_ _04076_ VPWR VGND _04100_ sg13g2_nor3_1
X_10372_ _01872_ _01681_ _04076_ VPWR VGND _04101_ sg13g2_nor3_1
X_10373_ _04100_ _04101_ _04061_ VPWR VGND _04102_ sg13g2_o21ai_1
X_10374_ _01877_ _04062_ VPWR VGND _04103_ sg13g2_nor2_1
X_10375_ _02491_ _04103_ _04101_ _04059_ VPWR VGND 
+ _04104_
+ sg13g2_a22oi_1
X_10376_ _04099_ _04102_ _04104_ VPWR VGND _04105_ sg13g2_nand3b_1
X_10377_ _01685_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[17]\ VPWR VGND _04106_ sg13g2_xor2_1
X_10378_ _04105_ _04106_ VPWR VGND _04107_ sg13g2_xnor2_1
X_10379_ _01897_ _04107_ VPWR VGND _04108_ sg13g2_xnor2_1
X_10380_ _02752_ _02278_ _04080_ VPWR VGND _04109_ sg13g2_mux2_1
X_10381_ _04108_ _04109_ VPWR VGND _04110_ sg13g2_nor2_1
X_10382_ _04070_ _04093_ _04110_ VPWR VGND _04111_ sg13g2_o21ai_1
X_10383_ _01895_ _04107_ VPWR VGND _04112_ sg13g2_or2_1
X_10384_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[17]\ VPWR VGND _04113_ sg13g2_inv_1
X_10385_ _01697_ _04113_ _04105_ VPWR VGND _04114_ sg13g2_a21oi_1
X_10386_ _02089_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[17]\ _04114_ VPWR VGND _04115_ sg13g2_a21oi_1
X_10387_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2081_o\ _04115_ _01902_ VPWR VGND _04116_ sg13g2_o21ai_1
X_10388_ _04111_ _04112_ _04116_ VPWR VGND _04117_ sg13g2_a21oi_1
X_10389_ _03949_ _03951_ _04117_ VPWR VGND _00457_ sg13g2_a21oi_1
X_10390_ _03947_ _02924_ VPWR VGND _04118_ sg13g2_nand2_1
X_10391_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2079_o[1]\ VPWR VGND _04119_ sg13g2_buf_1
X_10392_ _04119_ VPWR VGND _04120_ sg13g2_buf_1
X_10393_ _04120_ _01903_ VPWR VGND _04121_ sg13g2_nand2_1
X_10394_ _04118_ _04121_ _04117_ VPWR VGND _00458_ sg13g2_a21oi_1
X_10395_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[17]\ VPWR VGND _04122_ sg13g2_buf_1
X_10396_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[16]\ VPWR VGND _04123_ sg13g2_buf_1
X_10397_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[11]\ VPWR VGND _04124_ sg13g2_buf_1
X_10398_ _04124_ VPWR VGND _04125_ sg13g2_inv_1
X_10399_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[10]\ VPWR VGND _04126_ sg13g2_buf_1
X_10400_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[8]\ VPWR VGND _04127_ sg13g2_buf_1
X_10401_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[6]\ VPWR VGND _04128_ sg13g2_buf_1
X_10402_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[7]\ VPWR VGND _04129_ sg13g2_buf_1
X_10403_ _01609_ _04128_ _04129_ VPWR VGND _04130_ sg13g2_a21o_1
X_10404_ _01763_ _04129_ _04128_ VPWR VGND _04131_ sg13g2_and3_1
X_10405_ _01606_ _04127_ _04130_ _01614_ _04131_ VPWR 
+ VGND
+ _04132_ sg13g2_a221oi_1
X_10406_ _01606_ _04127_ VPWR VGND _04133_ sg13g2_nor2_1
X_10407_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[9]\ VPWR VGND _04134_ sg13g2_inv_1
X_10408_ _04132_ _04133_ _04134_ VPWR VGND _04135_ sg13g2_o21ai_1
X_10409_ _04134_ _04132_ _04133_ VPWR VGND _04136_ sg13g2_nor3_1
X_10410_ _01604_ _04135_ _04136_ VPWR VGND _04137_ sg13g2_a21o_1
X_10411_ _04126_ _04137_ VPWR VGND _04138_ sg13g2_nand2_1
X_10412_ _04126_ _04137_ _01648_ VPWR VGND _04139_ sg13g2_o21ai_1
X_10413_ _04139_ VPWR VGND _04140_ sg13g2_buf_1
X_10414_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[12]\ VPWR VGND _04141_ sg13g2_buf_1
X_10415_ _04141_ VPWR VGND _04142_ sg13g2_inv_1
X_10416_ _02018_ _04125_ _04138_ _04140_ _04142_ VPWR 
+ VGND
+ _04143_ sg13g2_a221oi_1
X_10417_ _02018_ _04142_ _04125_ VPWR VGND _04144_ sg13g2_nor3_1
X_10418_ _01661_ _04143_ _04144_ VPWR VGND _04145_ sg13g2_or3_1
X_10419_ _04145_ VPWR VGND _04146_ sg13g2_buf_1
X_10420_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[13]\ VPWR VGND _04147_ sg13g2_buf_1
X_10421_ _04147_ VPWR VGND _04148_ sg13g2_buf_1
X_10422_ _01639_ _04141_ VPWR VGND _04149_ sg13g2_nor2_1
X_10423_ _04138_ _04140_ _04149_ VPWR VGND _04150_ sg13g2_nand3_1
X_10424_ _04141_ _04124_ VPWR VGND _04151_ sg13g2_nor2_1
X_10425_ _04138_ _04140_ _04151_ VPWR VGND _04152_ sg13g2_nand3_1
X_10426_ _04125_ _04149_ VPWR VGND _04153_ sg13g2_nand2_1
X_10427_ _04148_ _04150_ _04152_ _04153_ VPWR VGND 
+ _04154_
+ sg13g2_and4_1
X_10428_ _04154_ VPWR VGND _04155_ sg13g2_buf_1
X_10429_ _04126_ VPWR VGND _04156_ sg13g2_inv_1
X_10430_ _01735_ _04135_ _04136_ VPWR VGND _04157_ sg13g2_a21oi_1
X_10431_ _04156_ _04157_ VPWR VGND _04158_ sg13g2_nand2_1
X_10432_ _04156_ _04157_ _01628_ VPWR VGND _04159_ sg13g2_o21ai_1
X_10433_ _04148_ _04141_ VPWR VGND _04160_ sg13g2_or2_1
X_10434_ _01661_ _04147_ VPWR VGND _04161_ sg13g2_or2_1
X_10435_ _04158_ _04159_ _04160_ _04161_ _04124_ VPWR 
+ VGND
+ _04162_ sg13g2_a221oi_1
X_10436_ _01639_ _04147_ VPWR VGND _04163_ sg13g2_nor2_1
X_10437_ _04142_ _04163_ VPWR VGND _04164_ sg13g2_nand2_1
X_10438_ _01661_ _01666_ VPWR VGND _04165_ sg13g2_nor2_1
X_10439_ _04148_ _04165_ VPWR VGND _04166_ sg13g2_nand2b_1
X_10440_ _04158_ _04159_ _04164_ _04166_ VPWR VGND 
+ _04167_
+ sg13g2_a22oi_1
X_10441_ _04148_ _04124_ VPWR VGND _04168_ sg13g2_nor2_1
X_10442_ _04151_ _04163_ _04168_ _04165_ VPWR VGND 
+ _04169_
+ sg13g2_a22oi_1
X_10443_ _04141_ _04161_ _04169_ VPWR VGND _04170_ sg13g2_o21ai_1
X_10444_ _01600_ _04162_ _04167_ _04170_ VPWR VGND 
+ _04171_
+ sg13g2_nor4_1
X_10445_ _04146_ _04155_ _04171_ VPWR VGND _04172_ sg13g2_a21o_1
X_10446_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[14]\ VPWR VGND _04173_ sg13g2_buf_1
X_10447_ _01672_ _04173_ VPWR VGND _04174_ sg13g2_or2_1
X_10448_ _04174_ VPWR VGND _04175_ sg13g2_buf_1
X_10449_ _01706_ _04173_ VPWR VGND _04176_ sg13g2_and2_1
X_10450_ _04172_ _04175_ _04176_ VPWR VGND _04177_ sg13g2_a21oi_1
X_10451_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[15]\ VPWR VGND _04178_ sg13g2_buf_1
X_10452_ _01876_ _04178_ VPWR VGND _04179_ sg13g2_nand2_1
X_10453_ _01876_ _04178_ VPWR VGND _04180_ sg13g2_nor2_1
X_10454_ _04177_ _04179_ _04180_ VPWR VGND _04181_ sg13g2_a21oi_1
X_10455_ _04123_ _04181_ _02343_ VPWR VGND _04182_ sg13g2_o21ai_1
X_10456_ _04123_ _04181_ VPWR VGND _04183_ sg13g2_nand2_1
X_10457_ _04182_ _04183_ VPWR VGND _04184_ sg13g2_nand2_1
X_10458_ _02089_ _04122_ _04184_ VPWR VGND _04185_ sg13g2_o21ai_1
X_10459_ _02089_ _04122_ VPWR VGND _04186_ sg13g2_nand2_1
X_10460_ _04185_ _04186_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2084_o\ VPWR VGND _04187_ sg13g2_a21oi_1
X_10461_ _01686_ _04122_ VPWR VGND _04188_ sg13g2_xor2_1
X_10462_ _04184_ _04188_ VPWR VGND _04189_ sg13g2_xnor2_1
X_10463_ _01681_ _04123_ VPWR VGND _04190_ sg13g2_xor2_1
X_10464_ _04181_ _04190_ VPWR VGND _04191_ sg13g2_xnor2_1
X_10465_ _04138_ _04140_ VPWR VGND _04192_ sg13g2_nand2_1
X_10466_ _01666_ _04124_ VPWR VGND _04193_ sg13g2_xnor2_1
X_10467_ _04192_ _04193_ VPWR VGND _04194_ sg13g2_xnor2_1
X_10468_ _01850_ _04194_ VPWR VGND _04195_ sg13g2_and2_1
X_10469_ _04195_ VPWR VGND _04196_ sg13g2_buf_1
X_10470_ _01730_ _04126_ VPWR VGND _04197_ sg13g2_xnor2_1
X_10471_ _04157_ _04197_ VPWR VGND _04198_ sg13g2_xnor2_1
X_10472_ _02197_ _04196_ _04198_ VPWR VGND _04199_ sg13g2_nor3_1
X_10473_ _02197_ _04198_ VPWR VGND _04200_ sg13g2_nand2_1
X_10474_ _04196_ _04200_ VPWR VGND _04201_ sg13g2_nor2_1
X_10475_ _04132_ _04133_ VPWR VGND _04202_ sg13g2_nor2_1
X_10476_ _01736_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[9]\ VPWR VGND _04203_ sg13g2_xor2_1
X_10477_ _04202_ _04203_ VPWR VGND _04204_ sg13g2_xnor2_1
X_10478_ _04204_ VPWR VGND _04205_ sg13g2_inv_1
X_10479_ _01959_ _04130_ _04131_ VPWR VGND _04206_ sg13g2_a21oi_1
X_10480_ _01990_ _04127_ VPWR VGND _04207_ sg13g2_xnor2_1
X_10481_ _04206_ _04207_ VPWR VGND _04208_ sg13g2_xnor2_1
X_10482_ _01754_ _04205_ _04208_ VPWR VGND _04209_ sg13g2_nor3_1
X_10483_ _02001_ _01754_ _04208_ VPWR VGND _04210_ sg13g2_nor3_1
X_10484_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[81]\ VPWR VGND _04211_ sg13g2_buf_1
X_10485_ _04211_ _02234_ _01983_ VPWR VGND _04212_ sg13g2_o21ai_1
X_10486_ _01818_ _04128_ VPWR VGND _04213_ sg13g2_xor2_1
X_10487_ _04211_ _02238_ _04213_ VPWR VGND _04214_ sg13g2_o21ai_1
X_10488_ _04212_ _04213_ _04214_ VPWR VGND _04215_ sg13g2_o21ai_1
X_10489_ _04215_ VPWR VGND _04216_ sg13g2_buf_1
X_10490_ _01792_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ VPWR VGND _04217_ sg13g2_nor2b_1
X_10491_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _04217_ _01797_ VPWR VGND _04218_ sg13g2_a21oi_1
X_10492_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _04217_ VPWR VGND _04219_ sg13g2_nor2_1
X_10493_ _01965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ VPWR VGND _04220_ sg13g2_nand2_1
X_10494_ _04218_ _04219_ _04220_ VPWR VGND _04221_ sg13g2_o21ai_1
X_10495_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ _01788_ VPWR VGND _04222_ sg13g2_nand2b_1
X_10496_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _04221_ _04222_ VPWR VGND 
+ _04223_
+ sg13g2_a22oi_1
X_10497_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _01783_ VPWR VGND _04224_ sg13g2_nand2b_1
X_10498_ _02222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _04224_ VPWR VGND _04225_ sg13g2_o21ai_1
X_10499_ _01809_ _04211_ VPWR VGND _04226_ sg13g2_nand2_1
X_10500_ _01809_ _04211_ VPWR VGND _04227_ sg13g2_or2_1
X_10501_ _04128_ _01773_ VPWR VGND _04228_ sg13g2_xor2_1
X_10502_ _01964_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _04226_ _04227_ _04228_ VPWR 
+ VGND
+ _04229_ sg13g2_a221oi_1
X_10503_ _04223_ _04225_ _04229_ VPWR VGND _04230_ sg13g2_o21ai_1
X_10504_ _04230_ VPWR VGND _04231_ sg13g2_buf_1
X_10505_ _01819_ _04128_ VPWR VGND _04232_ sg13g2_nand2_1
X_10506_ _01759_ _04129_ VPWR VGND _04233_ sg13g2_xor2_1
X_10507_ _04232_ _04233_ VPWR VGND _04234_ sg13g2_xnor2_1
X_10508_ _04216_ _04231_ _04234_ VPWR VGND _04235_ sg13g2_nand3_1
X_10509_ _04216_ _04231_ _04234_ VPWR VGND _04236_ sg13g2_a21oi_1
X_10510_ _02548_ _04235_ _04236_ VPWR VGND _04237_ sg13g2_a21o_1
X_10511_ _04209_ _04210_ _04237_ VPWR VGND _04238_ sg13g2_o21ai_1
X_10512_ _01814_ VPWR VGND _04239_ sg13g2_inv_1
X_10513_ _04239_ _04216_ _04231_ _04234_ VPWR VGND 
+ _04240_
+ sg13g2_nand4_1
X_10514_ _02548_ _01814_ VPWR VGND _04241_ sg13g2_nor2_1
X_10515_ _04216_ _04231_ _04241_ VPWR VGND _04242_ sg13g2_nand3_1
X_10516_ _04240_ _04242_ VPWR VGND _04243_ sg13g2_and2_1
X_10517_ _01989_ _04239_ _04234_ _04241_ VPWR VGND 
+ _04244_
+ sg13g2_a22oi_1
X_10518_ _04204_ _04208_ _04243_ _04244_ VPWR VGND 
+ _04245_
+ sg13g2_nand4_1
X_10519_ _02687_ _04208_ _04243_ _04244_ VPWR VGND 
+ _04246_
+ sg13g2_nand4_1
X_10520_ _02687_ _04204_ VPWR VGND _04247_ sg13g2_nand2_1
X_10521_ _04238_ _04245_ _04246_ _04247_ VPWR VGND 
+ _04248_
+ sg13g2_nand4_1
X_10522_ _04199_ _04201_ _04248_ VPWR VGND _04249_ sg13g2_o21ai_1
X_10523_ _02731_ _04194_ VPWR VGND _04250_ sg13g2_nor2_1
X_10524_ _04196_ _04198_ _02250_ VPWR VGND _04251_ sg13g2_nand3b_1
X_10525_ _04250_ _04251_ VPWR VGND _04252_ sg13g2_nor2b_1
X_10526_ _04138_ _04140_ _04125_ VPWR VGND _04253_ sg13g2_a21oi_1
X_10527_ _04125_ _04138_ _04140_ VPWR VGND _04254_ sg13g2_nand3_1
X_10528_ _01717_ _04253_ _04254_ VPWR VGND _04255_ sg13g2_o21ai_1
X_10529_ _01719_ _04141_ VPWR VGND _04256_ sg13g2_xor2_1
X_10530_ _04255_ _04256_ VPWR VGND _04257_ sg13g2_xnor2_1
X_10531_ _02571_ _04257_ VPWR VGND _04258_ sg13g2_nand2_1
X_10532_ _02571_ _04257_ VPWR VGND _04259_ sg13g2_or2_1
X_10533_ _04249_ _04252_ _04258_ _04259_ VPWR VGND 
+ _04260_
+ sg13g2_a22oi_1
X_10534_ _01719_ _04143_ _04144_ VPWR VGND _04261_ sg13g2_nor3_1
X_10535_ _04142_ _04255_ _04261_ VPWR VGND _04262_ sg13g2_a21oi_1
X_10536_ _01946_ _04148_ VPWR VGND _04263_ sg13g2_xor2_1
X_10537_ _04262_ _04263_ VPWR VGND _04264_ sg13g2_xnor2_1
X_10538_ _01913_ _04264_ VPWR VGND _04265_ sg13g2_nand2_1
X_10539_ _02572_ _04257_ _04265_ VPWR VGND _04266_ sg13g2_o21ai_1
X_10540_ _04148_ _04262_ VPWR VGND _04267_ sg13g2_nor2_1
X_10541_ _01912_ _01725_ _04267_ VPWR VGND _04268_ sg13g2_o21ai_1
X_10542_ _04173_ _01908_ VPWR VGND _04269_ sg13g2_xnor2_1
X_10543_ _04148_ _04150_ _04152_ _04153_ VPWR VGND 
+ _04270_
+ sg13g2_nand4_1
X_10544_ _04261_ _04270_ _02030_ VPWR VGND _04271_ sg13g2_o21ai_1
X_10545_ _04269_ _04271_ VPWR VGND _04272_ sg13g2_and2_1
X_10546_ _01658_ _04178_ VPWR VGND _04273_ sg13g2_xor2_1
X_10547_ _04177_ _04273_ VPWR VGND _04274_ sg13g2_xnor2_1
X_10548_ _02031_ _04146_ _04155_ VPWR VGND _04275_ sg13g2_nand3_1
X_10549_ _04172_ _04275_ _04269_ VPWR VGND _04276_ sg13g2_a21oi_1
X_10550_ _04268_ _04272_ _04274_ _02037_ _04276_ VPWR 
+ VGND
+ _04277_ sg13g2_a221oi_1
X_10551_ _04260_ _04266_ _04277_ VPWR VGND _04278_ sg13g2_o21ai_1
X_10552_ _01871_ _04173_ VPWR VGND _04279_ sg13g2_nor2_1
X_10553_ _04279_ _04176_ _02036_ VPWR VGND _04280_ sg13g2_o21ai_1
X_10554_ _01872_ _04173_ VPWR VGND _04281_ sg13g2_nand2_1
X_10555_ _04175_ _04281_ _04273_ VPWR VGND _04282_ sg13g2_nand3_1
X_10556_ _04146_ _04155_ _04171_ VPWR VGND _04283_ sg13g2_a21oi_1
X_10557_ _04280_ _04282_ _04283_ VPWR VGND _04284_ sg13g2_mux2_1
X_10558_ _02048_ _04283_ _01886_ VPWR VGND _04285_ sg13g2_o21ai_1
X_10559_ _04273_ _04285_ _04175_ VPWR VGND _04286_ sg13g2_nand3b_1
X_10560_ _04148_ _02630_ _03229_ VPWR VGND _04287_ sg13g2_a21o_1
X_10561_ _04279_ _04273_ VPWR VGND _04288_ sg13g2_and2_1
X_10562_ _04262_ _04287_ _04288_ VPWR VGND _04289_ sg13g2_o21ai_1
X_10563_ _03674_ _04270_ _04289_ VPWR VGND _04290_ sg13g2_a21oi_1
X_10564_ _02048_ _04289_ VPWR VGND _04291_ sg13g2_nand2_1
X_10565_ _02036_ _04290_ _04291_ VPWR VGND _04292_ sg13g2_o21ai_1
X_10566_ _04281_ _04273_ VPWR VGND _04293_ sg13g2_nor2_1
X_10567_ _01703_ _04172_ _04293_ VPWR VGND _04294_ sg13g2_o21ai_1
X_10568_ _04284_ _04286_ _04292_ _04294_ VPWR VGND 
+ _04295_
+ sg13g2_nand4_1
X_10569_ _01881_ _04191_ VPWR VGND _04296_ sg13g2_or2_1
X_10570_ _01881_ _04191_ VPWR VGND _04297_ sg13g2_nand2_1
X_10571_ _04278_ _04295_ _04296_ _04297_ VPWR VGND 
+ _04298_
+ sg13g2_a22oi_1
X_10572_ _02069_ _04191_ _04298_ VPWR VGND _04299_ sg13g2_a21o_1
X_10573_ _01897_ _04189_ VPWR VGND _04300_ sg13g2_xnor2_1
X_10574_ _02086_ _04189_ _04299_ _04300_ VPWR VGND 
+ _04301_
+ sg13g2_a22oi_1
X_10575_ _04187_ _04301_ _02108_ VPWR VGND _04302_ sg13g2_o21ai_1
X_10576_ _03950_ _02448_ VPWR VGND _04303_ sg13g2_nand2_1
X_10577_ _02099_ _04302_ _04303_ VPWR VGND _00459_ sg13g2_o21ai_1
X_10578_ _04120_ _02448_ VPWR VGND _04304_ sg13g2_nand2_1
X_10579_ _02106_ _04302_ _04304_ VPWR VGND _00460_ sg13g2_o21ai_1
X_10580_ _02103_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ sg13g2_buf_1
X_10581_ _01103_ _01693_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ VPWR VGND _00461_ sg13g2_a21oi_1
X_10582_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2099_o\ VPWR VGND _04305_ sg13g2_inv_1
X_10583_ _01104_ VPWR VGND _04306_ sg13g2_buf_1
X_10584_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2102_o\ _04306_ _02924_ VPWR VGND _04307_ sg13g2_nor3_1
X_10585_ _04305_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04307_ VPWR VGND _00462_ sg13g2_a21oi_1
X_10586_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2102_o\ VPWR VGND _04308_ sg13g2_inv_1
X_10587_ _02979_ _04306_ _02924_ VPWR VGND _04309_ sg13g2_nor3_1
X_10588_ _04308_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04309_ VPWR VGND _00463_ sg13g2_a21oi_1
X_10589_ _02979_ VPWR VGND _04310_ sg13g2_inv_1
X_10590_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2108_o\ _04306_ _02924_ VPWR VGND _04311_ sg13g2_nor3_1
X_10591_ _04310_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04311_ VPWR VGND _00464_ sg13g2_a21oi_1
X_10592_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2111_o\ _04306_ _02924_ VPWR VGND _04312_ sg13g2_nor3_1
X_10593_ _03241_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04312_ VPWR VGND _00465_ sg13g2_a21oi_1
X_10594_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2446_o\ _04306_ _02924_ VPWR VGND _04313_ sg13g2_nor3_1
X_10595_ _03307_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04313_ VPWR VGND _00466_ sg13g2_a21oi_1
X_10596_ _01104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2075_o\ _02924_ VPWR VGND _04314_ sg13g2_nor3_1
X_10597_ _01693_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04314_ VPWR VGND _00467_ sg13g2_a21oi_1
X_10598_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2075_o\ VPWR VGND _04315_ sg13g2_inv_1
X_10599_ _01104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2078_o\ _02924_ VPWR VGND _04316_ sg13g2_nor3_1
X_10600_ _04315_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04316_ VPWR VGND _00468_ sg13g2_a21oi_1
X_10601_ _01104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2081_o\ _02096_ VPWR VGND _04317_ sg13g2_nor3_1
X_10602_ _03790_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ _04317_ VPWR VGND _00469_ sg13g2_a21oi_1
X_10603_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2081_o\ VPWR VGND _04318_ sg13g2_inv_1
X_10604_ _02103_ VPWR VGND _04319_ sg13g2_buf_1
X_10605_ _01104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2084_o\ _02096_ VPWR VGND _04320_ sg13g2_nor3_1
X_10606_ _04318_ _04319_ _04320_ VPWR VGND _00470_ sg13g2_a21oi_1
X_10607_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2084_o\ VPWR VGND _04321_ sg13g2_inv_1
X_10608_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2087_o\ _04306_ _02096_ VPWR VGND _04322_ sg13g2_nor3_1
X_10609_ _04321_ _04319_ _04322_ VPWR VGND _00471_ sg13g2_a21oi_1
X_10610_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2087_o\ VPWR VGND _04323_ sg13g2_inv_1
X_10611_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2090_o\ _04306_ _02096_ VPWR VGND _04324_ sg13g2_nor3_1
X_10612_ _04323_ _04319_ _04324_ VPWR VGND _00472_ sg13g2_a21oi_1
X_10613_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2090_o\ VPWR VGND _04325_ sg13g2_inv_1
X_10614_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2093_o\ _04306_ _02096_ VPWR VGND _04326_ sg13g2_nor3_1
X_10615_ _04325_ _04319_ _04326_ VPWR VGND _00473_ sg13g2_a21oi_1
X_10616_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2096_o\ _04306_ _02096_ VPWR VGND _04327_ sg13g2_nor3_1
X_10617_ _02359_ _04319_ _04327_ VPWR VGND _00474_ sg13g2_a21oi_1
X_10618_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2096_o\ VPWR VGND _04328_ sg13g2_inv_1
X_10619_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2099_o\ _04306_ _02096_ VPWR VGND _04329_ sg13g2_nor3_1
X_10620_ _04328_ _04319_ _04329_ VPWR VGND _00475_ sg13g2_a21oi_1
X_10621_ \atbs_core_0.dac_control_0.dac_counter_value[0]\ VPWR VGND _04330_ sg13g2_buf_1
X_10622_ _00852_ _00951_ VPWR VGND _04331_ sg13g2_nand2_1
X_10623_ _01114_ _00858_ _00905_ VPWR VGND _04332_ sg13g2_a21oi_1
X_10624_ _04331_ _04332_ VPWR VGND _04333_ sg13g2_and2_1
X_10625_ _04333_ VPWR VGND _04334_ sg13g2_buf_1
X_10626_ _00047_ _04334_ VPWR VGND _04335_ sg13g2_nand2b_1
X_10627_ \atbs_core_0.dac_control_0.dac_counter_value[8]\ VPWR VGND _04336_ sg13g2_buf_2
X_10628_ _00037_ VPWR VGND _04337_ sg13g2_buf_2
X_10629_ _00041_ VPWR VGND _04338_ sg13g2_inv_1
X_10630_ _00855_ _01210_ VPWR VGND _04339_ sg13g2_nand2_1
X_10631_ _01321_ _01325_ _04339_ VPWR VGND _04340_ sg13g2_a21o_1
X_10632_ _04340_ VPWR VGND _04341_ sg13g2_buf_4
X_10633_ \atbs_core_0.debouncer_5.debounced\ \atbs_core_0.n1082_q\ _00853_ VPWR VGND _04342_ sg13g2_mux2_1
X_10634_ _04342_ VPWR VGND _04343_ sg13g2_buf_1
X_10635_ _00883_ _04343_ VPWR VGND _04344_ sg13g2_and2_1
X_10636_ _04344_ VPWR VGND _04345_ sg13g2_buf_1
X_10637_ \atbs_core_0.n1068_q[3]\ _04345_ VPWR VGND _04346_ sg13g2_nand2_1
X_10638_ _00855_ _01260_ _01317_ VPWR VGND _04347_ sg13g2_nand3_1
X_10639_ _04346_ _04347_ VPWR VGND _04348_ sg13g2_and2_1
X_10640_ _04348_ VPWR VGND _04349_ sg13g2_buf_1
X_10641_ _04338_ _04341_ _04349_ VPWR VGND _04350_ sg13g2_and3_1
X_10642_ _04350_ VPWR VGND _04351_ sg13g2_buf_2
X_10643_ _04341_ _04349_ _04338_ VPWR VGND _04352_ sg13g2_a21oi_1
X_10644_ _04351_ _04352_ VPWR VGND _04353_ sg13g2_nor2_2
X_10645_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ VPWR VGND _04354_ sg13g2_buf_1
X_10646_ \atbs_core_0.n1068_q[2]\ VPWR VGND _04355_ sg13g2_buf_1
X_10647_ _04355_ _04345_ VPWR VGND _04356_ sg13g2_nand2_1
X_10648_ _04356_ VPWR VGND _04357_ sg13g2_buf_1
X_10649_ _04354_ _04357_ VPWR VGND _04358_ sg13g2_nand2_1
X_10650_ _04354_ _00883_ VPWR VGND _04359_ sg13g2_nor2_1
X_10651_ _01210_ _01287_ _04359_ VPWR VGND _04360_ sg13g2_o21ai_1
X_10652_ _04358_ _04360_ _01302_ VPWR VGND _04361_ sg13g2_mux2_1
X_10653_ _04354_ _04357_ VPWR VGND _04362_ sg13g2_and2_1
X_10654_ _04354_ _00883_ _04357_ VPWR VGND _04363_ sg13g2_nand3_1
X_10655_ _04354_ _04357_ _04363_ VPWR VGND _04364_ sg13g2_o21ai_1
X_10656_ _01288_ _04362_ _04364_ VPWR VGND _04365_ sg13g2_a21oi_1
X_10657_ _04361_ _04365_ VPWR VGND _04366_ sg13g2_nand2_1
X_10658_ \atbs_core_0.n1068_q[1]\ _04345_ VPWR VGND _04367_ sg13g2_nand2_1
X_10659_ _04367_ VPWR VGND _04368_ sg13g2_buf_2
X_10660_ _00855_ _01253_ _01258_ _01263_ VPWR VGND 
+ _04369_
+ sg13g2_nand4_1
X_10661_ _04369_ VPWR VGND _04370_ sg13g2_buf_4
X_10662_ _00044_ VPWR VGND _04371_ sg13g2_buf_1
X_10663_ _04368_ _04370_ _04371_ VPWR VGND _04372_ sg13g2_a21oi_2
X_10664_ \atbs_core_0.dac_control_0.dac_counter_value[1]\ VPWR VGND _04373_ sg13g2_buf_1
X_10665_ _04373_ _04368_ VPWR VGND _04374_ sg13g2_nand2_1
X_10666_ _01253_ _01258_ _04374_ VPWR VGND _04375_ sg13g2_a21oi_1
X_10667_ _04373_ _00883_ VPWR VGND _04376_ sg13g2_nor2_1
X_10668_ _01253_ _01258_ _01263_ _04376_ VPWR VGND 
+ _04377_
+ sg13g2_and4_1
X_10669_ _01263_ _04374_ VPWR VGND _04378_ sg13g2_nor2_1
X_10670_ _04373_ _00883_ _04368_ VPWR VGND _04379_ sg13g2_nand3_1
X_10671_ _04373_ _04368_ _04379_ VPWR VGND _04380_ sg13g2_o21ai_1
X_10672_ _04375_ _04377_ _04378_ _04380_ VPWR VGND 
+ _04381_
+ sg13g2_or4_1
X_10673_ _00856_ _04343_ VPWR VGND _04382_ sg13g2_nor2_1
X_10674_ _04330_ _04382_ VPWR VGND _04383_ sg13g2_nand2_1
X_10675_ _04330_ _00856_ _01229_ _01232_ VPWR VGND 
+ _04384_
+ sg13g2_nand4_1
X_10676_ _01211_ _01224_ _04384_ VPWR VGND _04385_ sg13g2_a21o_1
X_10677_ _04361_ _04365_ _04383_ _04385_ VPWR VGND 
+ _04386_
+ sg13g2_a22oi_1
X_10678_ _01288_ _01302_ _00856_ VPWR VGND _04387_ sg13g2_nand3b_1
X_10679_ _00042_ VPWR VGND _04388_ sg13g2_buf_1
X_10680_ _04357_ _04387_ _04388_ VPWR VGND _04389_ sg13g2_a21oi_1
X_10681_ _04366_ _04372_ _04381_ _04386_ _04389_ VPWR 
+ VGND
+ _04390_ sg13g2_a221oi_1
X_10682_ _04390_ VPWR VGND _04391_ sg13g2_buf_2
X_10683_ _04341_ _04349_ VPWR VGND _04392_ sg13g2_nand2_1
X_10684_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ _04392_ VPWR VGND _04393_ sg13g2_nand2_1
X_10685_ _04353_ _04391_ _04393_ VPWR VGND _04394_ sg13g2_o21ai_1
X_10686_ _04394_ VPWR VGND _04395_ sg13g2_buf_4
X_10687_ \atbs_core_0.dac_control_0.dac_counter_value[4]\ VPWR VGND _04396_ sg13g2_buf_1
X_10688_ _04396_ VPWR VGND _04397_ sg13g2_inv_1
X_10689_ _04339_ VPWR VGND _04398_ sg13g2_inv_1
X_10690_ \atbs_core_0.n1068_q[4]\ _04345_ VPWR VGND _04399_ sg13g2_and2_1
X_10691_ _04399_ VPWR VGND _04400_ sg13g2_buf_1
X_10692_ _00856_ _01260_ _01344_ VPWR VGND _04401_ sg13g2_nand3_1
X_10693_ _04400_ _04401_ VPWR VGND _04402_ sg13g2_nand2b_1
X_10694_ _01351_ _04398_ _04402_ VPWR VGND _04403_ sg13g2_a21o_1
X_10695_ _04403_ VPWR VGND _04404_ sg13g2_buf_2
X_10696_ _04397_ _04404_ VPWR VGND _04405_ sg13g2_nor2_1
X_10697_ \atbs_core_0.n1068_q[5]\ _04345_ VPWR VGND _04406_ sg13g2_and2_1
X_10698_ _00856_ _01381_ _04406_ VPWR VGND _04407_ sg13g2_a21o_1
X_10699_ _01373_ _04398_ _04407_ VPWR VGND _04408_ sg13g2_a21o_1
X_10700_ _04408_ VPWR VGND _04409_ sg13g2_buf_2
X_10701_ _04337_ _04395_ _04405_ _04409_ VPWR VGND 
+ _04410_
+ sg13g2_nand4_1
X_10702_ _04337_ _04404_ _04409_ VPWR VGND _04411_ sg13g2_and3_1
X_10703_ _04351_ _04352_ _04397_ VPWR VGND _04412_ sg13g2_o21ai_1
X_10704_ _04396_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ VPWR VGND _04413_ sg13g2_nor2b_1
X_10705_ _00038_ VPWR VGND _04414_ sg13g2_inv_1
X_10706_ _04392_ _04413_ _04414_ VPWR VGND _04415_ sg13g2_a21oi_1
X_10707_ _04391_ _04412_ _04415_ VPWR VGND _04416_ sg13g2_o21ai_1
X_10708_ \atbs_core_0.dac_control_0.dac_counter_value[5]\ _04409_ _04411_ _04416_ VPWR VGND 
+ _04417_
+ sg13g2_a22oi_1
X_10709_ _04337_ _04409_ VPWR VGND _04418_ sg13g2_nor2_1
X_10710_ _04404_ _04418_ VPWR VGND _04419_ sg13g2_and2_1
X_10711_ _04405_ _04418_ VPWR VGND _04420_ sg13g2_and2_1
X_10712_ _04416_ _04419_ _04420_ _04395_ VPWR VGND 
+ _04421_
+ sg13g2_a22oi_1
X_10713_ \atbs_core_0.dac_control_0.dac_counter_value[7]\ VPWR VGND _04422_ sg13g2_buf_1
X_10714_ _00944_ _01430_ VPWR VGND _04423_ sg13g2_nor2_1
X_10715_ _04423_ VPWR VGND _04424_ sg13g2_buf_1
X_10716_ _00858_ _01407_ VPWR VGND _04425_ sg13g2_and2_1
X_10717_ _04425_ VPWR VGND _04426_ sg13g2_buf_1
X_10718_ _04422_ _04424_ _04426_ VPWR VGND _04427_ sg13g2_a21oi_1
X_10719_ _04410_ _04417_ _04421_ _04427_ VPWR VGND 
+ _04428_
+ sg13g2_nand4_1
X_10720_ \atbs_core_0.dac_control_0.dac_counter_value[6]\ VPWR VGND _04429_ sg13g2_buf_1
X_10721_ \atbs_core_0.dac_control_0.dac_counter_value[7]\ _04424_ _04429_ VPWR VGND _04430_ sg13g2_a21oi_1
X_10722_ _04410_ _04417_ _04421_ _04430_ VPWR VGND 
+ _04431_
+ sg13g2_nand4_1
X_10723_ _04422_ _04424_ VPWR VGND _04432_ sg13g2_nand2_1
X_10724_ _04429_ VPWR VGND _04433_ sg13g2_buf_1
X_10725_ _04433_ _04426_ VPWR VGND _04434_ sg13g2_nor2_1
X_10726_ _04422_ _04424_ VPWR VGND _04435_ sg13g2_nor2_1
X_10727_ _04432_ _04434_ _04435_ VPWR VGND _04436_ sg13g2_a21oi_1
X_10728_ _04428_ _04431_ _04436_ VPWR VGND _04437_ sg13g2_and3_2
X_10729_ _04437_ VPWR VGND _04438_ sg13g2_buf_4
X_10730_ _04336_ _04438_ VPWR VGND _04439_ sg13g2_xnor2_1
X_10731_ _00823_ _00852_ _00951_ VPWR VGND _04440_ sg13g2_nand3_1
X_10732_ _04335_ _04439_ _04440_ VPWR VGND _04441_ sg13g2_o21ai_1
X_10733_ _04441_ VPWR VGND _04442_ sg13g2_buf_4
X_10734_ _04442_ VPWR VGND _04443_ sg13g2_buf_8
X_10735_ _00824_ VPWR VGND _04444_ sg13g2_buf_2
X_10736_ _04334_ VPWR VGND _04445_ sg13g2_buf_1
X_10737_ _00858_ _01235_ _04382_ VPWR VGND _04446_ sg13g2_a21oi_1
X_10738_ _04330_ _04446_ VPWR VGND _04447_ sg13g2_xnor2_1
X_10739_ _04422_ VPWR VGND _04448_ sg13g2_inv_1
X_10740_ _00857_ _01400_ _01405_ VPWR VGND _04449_ sg13g2_nand3_1
X_10741_ _04449_ VPWR VGND _04450_ sg13g2_buf_1
X_10742_ _04429_ _04450_ VPWR VGND _04451_ sg13g2_xnor2_1
X_10743_ _00857_ _01303_ _04345_ _04355_ _04388_ VPWR 
+ VGND
+ _04452_ sg13g2_a221oi_1
X_10744_ _04355_ _04345_ VPWR VGND _04453_ sg13g2_and2_1
X_10745_ _04453_ VPWR VGND _04454_ sg13g2_buf_1
X_10746_ _01283_ _01286_ VPWR VGND _04455_ sg13g2_xor2_1
X_10747_ _04388_ _00857_ VPWR VGND _04456_ sg13g2_nand2_1
X_10748_ _01260_ _04455_ _04456_ VPWR VGND _04457_ sg13g2_a21oi_1
X_10749_ _04388_ _04454_ _04457_ _01302_ VPWR VGND 
+ _04458_
+ sg13g2_a22oi_1
X_10750_ _04452_ _04458_ VPWR VGND _04459_ sg13g2_nand2b_1
X_10751_ _04371_ _04368_ _04370_ VPWR VGND _04460_ sg13g2_and3_1
X_10752_ _04372_ _04460_ VPWR VGND _04461_ sg13g2_nor2_1
X_10753_ _04336_ _04451_ _04459_ _04461_ VPWR VGND 
+ _04462_
+ sg13g2_nor4_1
X_10754_ _04337_ _04409_ VPWR VGND _04463_ sg13g2_xor2_1
X_10755_ _00069_ _04446_ VPWR VGND _04464_ sg13g2_xnor2_1
X_10756_ _04414_ _04404_ VPWR VGND _04465_ sg13g2_xnor2_1
X_10757_ _04353_ _04463_ _04464_ _04465_ VPWR VGND 
+ _04466_
+ sg13g2_and4_1
X_10758_ _04337_ _04409_ VPWR VGND _04467_ sg13g2_nand2_1
X_10759_ _04433_ _04467_ VPWR VGND _04468_ sg13g2_nand2_1
X_10760_ _04462_ _04466_ _04468_ VPWR VGND _04469_ sg13g2_a21oi_1
X_10761_ _04337_ _04409_ _04462_ _04466_ _04426_ VPWR 
+ VGND
+ _04470_ sg13g2_a221oi_1
X_10762_ _04368_ _04370_ VPWR VGND _04471_ sg13g2_nand2_1
X_10763_ _00069_ _00856_ VPWR VGND _04472_ sg13g2_nand2_1
X_10764_ _01224_ _01233_ _04472_ VPWR VGND _04473_ sg13g2_or3_1
X_10765_ _04473_ VPWR VGND _04474_ sg13g2_buf_1
X_10766_ _01219_ _01227_ _01228_ VPWR VGND _04475_ sg13g2_a21o_1
X_10767_ _01211_ _04475_ _01231_ _04472_ VPWR VGND 
+ _04476_
+ sg13g2_nor4_1
X_10768_ _00069_ _04382_ _04476_ VPWR VGND _04477_ sg13g2_a21oi_1
X_10769_ _04371_ VPWR VGND _04478_ sg13g2_inv_1
X_10770_ _04474_ _04477_ _04478_ VPWR VGND _04479_ sg13g2_a21oi_1
X_10771_ _04478_ _04474_ _04477_ VPWR VGND _04480_ sg13g2_nand3_1
X_10772_ _04471_ _04479_ _04480_ VPWR VGND _04481_ sg13g2_o21ai_1
X_10773_ _00038_ _04392_ VPWR VGND _04482_ sg13g2_nand2_1
X_10774_ _00038_ _00041_ VPWR VGND _04483_ sg13g2_nand2_1
X_10775_ _04458_ _04481_ _04482_ _04483_ _04452_ VPWR 
+ VGND
+ _04484_ sg13g2_a221oi_1
X_10776_ _04357_ _04387_ VPWR VGND _04485_ sg13g2_nand2_1
X_10777_ _04474_ _04477_ VPWR VGND _04486_ sg13g2_nand2_1
X_10778_ _04388_ _04485_ _04486_ _04371_ _04471_ VPWR 
+ VGND
+ _04487_ sg13g2_a221oi_1
X_10779_ _04487_ VPWR VGND _04488_ sg13g2_buf_1
X_10780_ _04478_ _04458_ _04474_ _04477_ VPWR VGND 
+ _04489_
+ sg13g2_nand4_1
X_10781_ _04452_ _04489_ VPWR VGND _04490_ sg13g2_nand2b_1
X_10782_ _04404_ _04392_ VPWR VGND _04491_ sg13g2_nand2_1
X_10783_ _04488_ _04490_ _04491_ VPWR VGND _04492_ sg13g2_nor3_1
X_10784_ _00041_ _04404_ VPWR VGND _04493_ sg13g2_nand2_1
X_10785_ _04488_ _04490_ _04493_ VPWR VGND _04494_ sg13g2_nor3_1
X_10786_ _04341_ _04349_ _04483_ VPWR VGND _04495_ sg13g2_a21oi_1
X_10787_ _00038_ _04404_ _04495_ VPWR VGND _04496_ sg13g2_a21oi_1
X_10788_ _04338_ _04491_ _04496_ VPWR VGND _04497_ sg13g2_o21ai_1
X_10789_ _04484_ _04492_ _04494_ _04497_ VPWR VGND 
+ _04498_
+ sg13g2_nor4_2
X_10790_ _04469_ _04470_ _04498_ VPWR VGND _04499_ sg13g2_o21ai_1
X_10791_ _04433_ _04450_ VPWR VGND _04500_ sg13g2_nand2_1
X_10792_ _04433_ _04450_ _04418_ VPWR VGND _04501_ sg13g2_o21ai_1
X_10793_ _04500_ _04501_ VPWR VGND _04502_ sg13g2_and2_1
X_10794_ _04448_ _04424_ _04499_ _04502_ VPWR VGND 
+ _04503_
+ sg13g2_a22oi_1
X_10795_ _04337_ _04409_ VPWR VGND _04504_ sg13g2_xnor2_1
X_10796_ _04336_ VPWR VGND _04505_ sg13g2_inv_1
X_10797_ _04372_ _04460_ _04505_ VPWR VGND _04506_ sg13g2_o21ai_1
X_10798_ _04504_ _04451_ _04459_ _04506_ VPWR VGND 
+ _04507_
+ sg13g2_or4_1
X_10799_ _04353_ _04464_ _04465_ VPWR VGND _04508_ sg13g2_nand3_1
X_10800_ _00070_ VPWR VGND _04509_ sg13g2_inv_1
X_10801_ _04507_ _04508_ _04509_ VPWR VGND _04510_ sg13g2_o21ai_1
X_10802_ _00944_ _01430_ VPWR VGND _04511_ sg13g2_or2_1
X_10803_ _04511_ VPWR VGND _04512_ sg13g2_buf_1
X_10804_ _04422_ _00070_ _04512_ VPWR VGND _04513_ sg13g2_nor3_1
X_10805_ _04422_ _04512_ _04513_ VPWR VGND _04514_ sg13g2_a21oi_1
X_10806_ _04510_ _04514_ VPWR VGND _04515_ sg13g2_nand2_1
X_10807_ _04503_ _04515_ VPWR VGND _04516_ sg13g2_or2_1
X_10808_ _04516_ VPWR VGND _04517_ sg13g2_buf_1
X_10809_ _04445_ _04464_ VPWR VGND _04518_ sg13g2_nor2_1
X_10810_ _04445_ _04447_ _04517_ _04518_ VPWR VGND 
+ _04519_
+ sg13g2_a22oi_1
X_10811_ _04444_ _04442_ _04519_ VPWR VGND _04520_ sg13g2_nor3_1
X_10812_ _04330_ _04443_ _04520_ VPWR VGND _00484_ sg13g2_a21o_1
X_10813_ _04499_ _04502_ VPWR VGND _04521_ sg13g2_nand2_1
X_10814_ _04521_ VPWR VGND _04522_ sg13g2_buf_2
X_10815_ _04448_ _04424_ _04334_ VPWR VGND _04523_ sg13g2_a21oi_1
X_10816_ _04478_ _04486_ VPWR VGND _04524_ sg13g2_xnor2_1
X_10817_ _04510_ _04514_ _04334_ VPWR VGND _04525_ sg13g2_a21o_1
X_10818_ _04525_ VPWR VGND _04526_ sg13g2_buf_1
X_10819_ _04383_ _04385_ VPWR VGND _04527_ sg13g2_nand2_1
X_10820_ _04373_ _04527_ VPWR VGND _04528_ sg13g2_xor2_1
X_10821_ _04334_ _04528_ _04471_ VPWR VGND _04529_ sg13g2_a21oi_1
X_10822_ _04524_ _04526_ _04529_ VPWR VGND _04530_ sg13g2_o21ai_1
X_10823_ _04331_ _04332_ VPWR VGND _04531_ sg13g2_nand2_1
X_10824_ _04531_ _04528_ _04471_ VPWR VGND _04532_ sg13g2_o21ai_1
X_10825_ _04532_ _04526_ VPWR VGND _04533_ sg13g2_nand2b_1
X_10826_ _04522_ _04523_ _04530_ _04533_ VPWR VGND 
+ _04534_
+ sg13g2_a22oi_1
X_10827_ _04524_ _04529_ VPWR VGND _04535_ sg13g2_nand2_1
X_10828_ _04524_ _04532_ _04535_ VPWR VGND _04536_ sg13g2_o21ai_1
X_10829_ _04444_ _04534_ _04536_ VPWR VGND _04537_ sg13g2_nor3_1
X_10830_ _04444_ \atbs_core_0.dac_control_0.dac_init_value[1]\ _04537_ VPWR VGND _04538_ sg13g2_a21oi_1
X_10831_ _04373_ _04443_ VPWR VGND _04539_ sg13g2_nand2_1
X_10832_ _04443_ _04538_ _04539_ VPWR VGND _00485_ sg13g2_o21ai_1
X_10833_ _04481_ _04459_ VPWR VGND _04540_ sg13g2_xor2_1
X_10834_ _04445_ _04540_ VPWR VGND _04541_ sg13g2_nor2_1
X_10835_ _04527_ _04381_ _04372_ VPWR VGND _04542_ sg13g2_a21o_1
X_10836_ _04366_ _04542_ VPWR VGND _04543_ sg13g2_xor2_1
X_10837_ _04517_ _04541_ _04543_ _04445_ VPWR VGND 
+ _04544_
+ sg13g2_a22oi_1
X_10838_ _00823_ \atbs_core_0.dac_control_0.dac_init_value[2]\ VPWR VGND _04545_ sg13g2_nor2_1
X_10839_ _00823_ _04544_ _04545_ VPWR VGND _04546_ sg13g2_a21oi_1
X_10840_ _04546_ _04354_ _04443_ VPWR VGND _00486_ sg13g2_mux2_1
X_10841_ \atbs_core_0.dac_control_0.dac_init_value[3]\ VPWR VGND _04547_ sg13g2_inv_1
X_10842_ _04488_ _04490_ VPWR VGND _04548_ sg13g2_nor2_1
X_10843_ _04548_ _04522_ _04523_ VPWR VGND _04549_ sg13g2_and3_1
X_10844_ _04391_ _04334_ VPWR VGND _04550_ sg13g2_nand2b_1
X_10845_ _04353_ _04550_ VPWR VGND _04551_ sg13g2_and2_1
X_10846_ _04531_ _04548_ _04515_ VPWR VGND _04552_ sg13g2_nand3_1
X_10847_ _04551_ _04552_ VPWR VGND _04553_ sg13g2_nand2_1
X_10848_ _04445_ _04391_ _04353_ VPWR VGND _04554_ sg13g2_a21oi_1
X_10849_ _04548_ _04526_ _04554_ VPWR VGND _04555_ sg13g2_o21ai_1
X_10850_ _04549_ _04553_ _04555_ VPWR VGND _04556_ sg13g2_o21ai_1
X_10851_ _04548_ _04551_ VPWR VGND _04557_ sg13g2_nor2_1
X_10852_ _04522_ _04523_ _04557_ VPWR VGND _04558_ sg13g2_nand3_1
X_10853_ _00823_ _04558_ VPWR VGND _04559_ sg13g2_and2_1
X_10854_ _04444_ _04547_ _04556_ _04559_ _04442_ VPWR 
+ VGND
+ _04560_ sg13g2_a221oi_1
X_10855_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ _04443_ _04560_ VPWR VGND _00487_ sg13g2_a21o_1
X_10856_ _04352_ _04548_ VPWR VGND _04561_ sg13g2_nor2_1
X_10857_ _04351_ _04561_ VPWR VGND _04562_ sg13g2_nor2_1
X_10858_ _04562_ _04465_ VPWR VGND _04563_ sg13g2_xor2_1
X_10859_ _04445_ _04563_ VPWR VGND _04564_ sg13g2_nor2_1
X_10860_ _04396_ _04404_ VPWR VGND _04565_ sg13g2_xnor2_1
X_10861_ _04395_ _04565_ VPWR VGND _04566_ sg13g2_xnor2_1
X_10862_ _04517_ _04564_ _04566_ _04445_ VPWR VGND 
+ _04567_
+ sg13g2_a22oi_1
X_10863_ _00823_ \atbs_core_0.dac_control_0.dac_init_value[4]\ VPWR VGND _04568_ sg13g2_nor2_1
X_10864_ _00823_ _04567_ _04568_ VPWR VGND _04569_ sg13g2_a21oi_1
X_10865_ _04569_ _04396_ _04443_ VPWR VGND _00488_ sg13g2_mux2_1
X_10866_ \atbs_core_0.dac_control_0.dac_counter_value[5]\ VPWR VGND _04570_ sg13g2_inv_1
X_10867_ _04404_ _04416_ _04405_ _04395_ VPWR VGND 
+ _04571_
+ sg13g2_a22oi_1
X_10868_ _04445_ _04571_ VPWR VGND _04572_ sg13g2_nand2_1
X_10869_ _04484_ _04492_ _04494_ _04497_ VPWR VGND 
+ _04573_
+ sg13g2_or4_1
X_10870_ _04573_ _04526_ VPWR VGND _04574_ sg13g2_or2_1
X_10871_ _04504_ _04572_ _04574_ VPWR VGND _04575_ sg13g2_nand3_1
X_10872_ _04498_ _04522_ _04523_ VPWR VGND _04576_ sg13g2_and3_1
X_10873_ _04531_ _04571_ VPWR VGND _04577_ sg13g2_nor2_1
X_10874_ _04498_ _04526_ _04463_ VPWR VGND _04578_ sg13g2_o21ai_1
X_10875_ _04577_ _04578_ VPWR VGND _04579_ sg13g2_or2_1
X_10876_ _04575_ _04576_ _04579_ VPWR VGND _04580_ sg13g2_o21ai_1
X_10877_ _04573_ _04522_ _04523_ _04575_ VPWR VGND 
+ _04581_
+ sg13g2_nand4_1
X_10878_ _04580_ _04581_ _04444_ VPWR VGND _04582_ sg13g2_a21o_1
X_10879_ _04444_ \atbs_core_0.dac_control_0.dac_init_value[5]\ _04443_ VPWR VGND _04583_ sg13g2_a21oi_1
X_10880_ _04570_ _04443_ _04582_ _04583_ VPWR VGND 
+ _00489_
+ sg13g2_a22oi_1
X_10881_ _04410_ _04417_ _04421_ VPWR VGND _04584_ sg13g2_nand3_1
X_10882_ _04584_ VPWR VGND _04585_ sg13g2_buf_1
X_10883_ _04585_ _04451_ VPWR VGND _04586_ sg13g2_xor2_1
X_10884_ _00824_ _04531_ VPWR VGND _04587_ sg13g2_nor2_1
X_10885_ _04418_ _04498_ _04467_ VPWR VGND _04588_ sg13g2_o21ai_1
X_10886_ _04426_ _04588_ VPWR VGND _04589_ sg13g2_xnor2_1
X_10887_ _00824_ _04445_ VPWR VGND _04590_ sg13g2_nor2_1
X_10888_ _04503_ _04515_ _04590_ VPWR VGND _04591_ sg13g2_o21ai_1
X_10889_ _04591_ VPWR VGND _04592_ sg13g2_buf_1
X_10890_ _04433_ _04589_ _04592_ VPWR VGND _04593_ sg13g2_nor3_1
X_10891_ _04444_ \atbs_core_0.dac_control_0.dac_init_value[6]\ _04586_ _04587_ _04593_ VPWR 
+ VGND
+ _04594_ sg13g2_a221oi_1
X_10892_ _04433_ _04589_ VPWR VGND _04595_ sg13g2_nand2_1
X_10893_ _04592_ _04595_ VPWR VGND _04596_ sg13g2_nor2_1
X_10894_ _04433_ _04442_ _04596_ VPWR VGND _04597_ sg13g2_a21oi_1
X_10895_ _04443_ _04594_ _04597_ VPWR VGND _00490_ sg13g2_o21ai_1
X_10896_ _04426_ _04585_ _04433_ VPWR VGND _04598_ sg13g2_a21o_1
X_10897_ _04426_ _04585_ _04598_ VPWR VGND _04599_ sg13g2_o21ai_1
X_10898_ _04448_ _04424_ VPWR VGND _04600_ sg13g2_xnor2_1
X_10899_ _04599_ _04600_ VPWR VGND _04601_ sg13g2_xnor2_1
X_10900_ _04433_ _04450_ VPWR VGND _04602_ sg13g2_nor2_1
X_10901_ _04500_ _04588_ _04602_ VPWR VGND _04603_ sg13g2_a21oi_1
X_10902_ _04512_ _04603_ VPWR VGND _04604_ sg13g2_xnor2_1
X_10903_ _04422_ _04592_ _04604_ VPWR VGND _04605_ sg13g2_nor3_1
X_10904_ _04444_ \atbs_core_0.dac_control_0.dac_init_value[7]\ _04587_ _04601_ _04605_ VPWR 
+ VGND
+ _04606_ sg13g2_a221oi_1
X_10905_ _04592_ _04604_ VPWR VGND _04607_ sg13g2_nor2b_1
X_10906_ _04442_ _04607_ _04422_ VPWR VGND _04608_ sg13g2_o21ai_1
X_10907_ _04443_ _04606_ _04608_ VPWR VGND _00491_ sg13g2_o21ai_1
X_10908_ _04336_ _04335_ VPWR VGND _04609_ sg13g2_nor2_1
X_10909_ _04438_ _04609_ VPWR VGND _04610_ sg13g2_and2_1
X_10910_ _04335_ _04438_ _04440_ VPWR VGND _04611_ sg13g2_o21ai_1
X_10911_ _04444_ \atbs_core_0.dac_control_0.dac_init_value[8]\ _04611_ _04336_ VPWR VGND 
+ _04612_
+ sg13g2_a22oi_1
X_10912_ _04512_ _04522_ VPWR VGND _04613_ sg13g2_nor2_1
X_10913_ _04512_ _04522_ _04422_ VPWR VGND _04614_ sg13g2_a21oi_1
X_10914_ _00070_ _04445_ _04613_ _04614_ VPWR VGND 
+ _04615_
+ sg13g2_nor4_1
X_10915_ _04531_ _04439_ VPWR VGND _04616_ sg13g2_nor2_1
X_10916_ _00852_ _00951_ _04438_ _04609_ _04444_ VPWR 
+ VGND
+ _04617_ sg13g2_a221oi_1
X_10917_ _04615_ _04616_ _04617_ VPWR VGND _04618_ sg13g2_o21ai_1
X_10918_ _04610_ _04612_ _04618_ VPWR VGND _00492_ sg13g2_o21ai_1
X_10919_ \atbs_core_0.dac_control_0.dac_wr_o\ VPWR VGND _04619_ sg13g2_buf_1
X_10920_ dac_upper_o[0] _04330_ _04619_ VPWR VGND _00493_ sg13g2_mux2_1
X_10921_ dac_upper_o[1] _04373_ _04619_ VPWR VGND _00494_ sg13g2_mux2_1
X_10922_ dac_upper_o[2] _04354_ _04619_ VPWR VGND _00495_ sg13g2_mux2_1
X_10923_ dac_upper_o[3] \atbs_core_0.dac_control_0.dac_counter_value[3]\ _04619_ VPWR VGND _00496_ sg13g2_mux2_1
X_10924_ dac_upper_o[4] _04396_ _04619_ VPWR VGND _00497_ sg13g2_mux2_1
X_10925_ dac_upper_o[5] \atbs_core_0.dac_control_0.dac_counter_value[5]\ _04619_ VPWR VGND _00498_ sg13g2_mux2_1
X_10926_ dac_upper_o[6] _04433_ _04619_ VPWR VGND _00499_ sg13g2_mux2_1
X_10927_ dac_upper_o[7] _04422_ _04619_ VPWR VGND _00500_ sg13g2_mux2_1
X_10928_ \atbs_core_0.dac_control_0.n1592_q[1]\ \atbs_core_0.dac_control_0.n1592_q[0]\ VPWR VGND _04620_ sg13g2_nand2_1
X_10929_ _00030_ _04620_ VPWR VGND _04621_ sg13g2_or2_1
X_10930_ \atbs_core_0.dac_control_0.dac_change_in_progress\ _04621_ \atbs_core_0.dac_control_0.dac_counter_strb\ VPWR VGND _00501_ sg13g2_a21o_1
X_10931_ \atbs_core_0.dac_control_1.dac_counter_value[8]\ VPWR VGND _04622_ sg13g2_inv_1
X_10932_ \atbs_core_0.dac_control_1.dac_counter_value[7]\ VPWR VGND _04623_ sg13g2_buf_1
X_10933_ _00944_ _01555_ VPWR VGND _04624_ sg13g2_nor2_1
X_10934_ _04623_ _04624_ VPWR VGND _04625_ sg13g2_nor2_1
X_10935_ _04623_ _04624_ VPWR VGND _04626_ sg13g2_and2_1
X_10936_ _01023_ _01206_ _01321_ _01325_ _00944_ VPWR 
+ VGND
+ _04627_ sg13g2_a221oi_1
X_10937_ _00856_ _01317_ VPWR VGND _04628_ sg13g2_nand2_1
X_10938_ _01498_ _04628_ _04346_ VPWR VGND _04629_ sg13g2_o21ai_1
X_10939_ _04627_ _04629_ VPWR VGND _04630_ sg13g2_nor2_1
X_10940_ _04630_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ VPWR VGND _04631_ sg13g2_nor2b_1
X_10941_ \atbs_core_0.dac_control_1.dac_counter_value[0]\ VPWR VGND _04632_ sg13g2_buf_4
X_10942_ \atbs_core_0.dac_control_1.dac_counter_value[2]\ VPWR VGND _04633_ sg13g2_buf_1
X_10943_ _04633_ _04357_ VPWR VGND _04634_ sg13g2_and2_1
X_10944_ _01484_ _01498_ _04634_ VPWR VGND _04635_ sg13g2_nand3_1
X_10945_ _04633_ _00883_ _04455_ _01449_ VPWR VGND 
+ _04636_
+ sg13g2_nor4_1
X_10946_ _01485_ _04634_ _04636_ VPWR VGND _04637_ sg13g2_a21oi_1
X_10947_ _04633_ _00944_ VPWR VGND _04638_ sg13g2_nand2_1
X_10948_ _04633_ _04638_ _04357_ VPWR VGND _04639_ sg13g2_mux2_1
X_10949_ _04633_ _00944_ _01484_ _01485_ VPWR VGND 
+ _04640_
+ sg13g2_or4_1
X_10950_ _04635_ _04637_ _04639_ _04640_ VPWR VGND 
+ _04641_
+ sg13g2_nand4_1
X_10951_ \atbs_core_0.n1068_q[1]\ _04345_ VPWR VGND _04642_ sg13g2_and2_1
X_10952_ _01462_ _01463_ _01465_ _04642_ VPWR VGND 
+ _04643_
+ sg13g2_nor4_1
X_10953_ _01262_ _01462_ _04368_ VPWR VGND _04644_ sg13g2_and3_1
X_10954_ _00883_ _04368_ _04643_ _01468_ _04644_ VPWR 
+ VGND
+ _04645_ sg13g2_a221oi_1
X_10955_ _04645_ VPWR VGND _04646_ sg13g2_buf_2
X_10956_ \atbs_core_0.dac_control_1.dac_counter_value[1]\ _04646_ VPWR VGND _04647_ sg13g2_xor2_1
X_10957_ _00856_ _01453_ _04382_ VPWR VGND _04648_ sg13g2_a21o_1
X_10958_ _04648_ VPWR VGND _04649_ sg13g2_buf_4
X_10959_ _04632_ _04641_ _04647_ _04649_ VPWR VGND 
+ _04650_
+ sg13g2_nand4_1
X_10960_ _00058_ VPWR VGND _04651_ sg13g2_inv_1
X_10961_ _00857_ _01487_ _04454_ VPWR VGND _04652_ sg13g2_a21o_1
X_10962_ _00059_ VPWR VGND _04653_ sg13g2_inv_1
X_10963_ _04653_ _04646_ VPWR VGND _04654_ sg13g2_and2_1
X_10964_ _04651_ _04652_ _04641_ _04654_ VPWR VGND 
+ _04655_
+ sg13g2_a22oi_1
X_10965_ _04627_ _04629_ _00057_ VPWR VGND _04656_ sg13g2_o21ai_1
X_10966_ _04656_ VPWR VGND _04657_ sg13g2_buf_1
X_10967_ _00057_ VPWR VGND _04658_ sg13g2_inv_1
X_10968_ _04658_ _04630_ VPWR VGND _04659_ sg13g2_nand2_1
X_10969_ _04650_ _04655_ _04657_ _04659_ VPWR VGND 
+ _04660_
+ sg13g2_a22oi_1
X_10970_ \atbs_core_0.dac_control_1.dac_counter_value[4]\ VPWR VGND _04661_ sg13g2_buf_1
X_10971_ _04661_ VPWR VGND _04662_ sg13g2_inv_1
X_10972_ _00857_ _01514_ _04400_ VPWR VGND _04663_ sg13g2_a21o_1
X_10973_ _04663_ VPWR VGND _04664_ sg13g2_buf_2
X_10974_ _04662_ _04664_ VPWR VGND _04665_ sg13g2_nor2_1
X_10975_ _04631_ _04660_ _04665_ VPWR VGND _04666_ sg13g2_o21ai_1
X_10976_ _04666_ VPWR VGND _04667_ sg13g2_buf_2
X_10977_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ _04662_ VPWR VGND _04668_ sg13g2_nand2_1
X_10978_ _00056_ VPWR VGND _04669_ sg13g2_buf_1
X_10979_ _04630_ _04668_ _04669_ VPWR VGND _04670_ sg13g2_o21ai_1
X_10980_ _04650_ _04655_ _04657_ _04659_ _04661_ VPWR 
+ VGND
+ _04671_ sg13g2_a221oi_1
X_10981_ _04670_ _04671_ _04664_ VPWR VGND _04672_ sg13g2_o21ai_1
X_10982_ _04672_ VPWR VGND _04673_ sg13g2_buf_4
X_10983_ _00055_ VPWR VGND _04674_ sg13g2_buf_1
X_10984_ _00858_ _01524_ _04406_ VPWR VGND _04675_ sg13g2_a21o_1
X_10985_ _04675_ VPWR VGND _04676_ sg13g2_buf_1
X_10986_ _04676_ VPWR VGND _04677_ sg13g2_buf_1
X_10987_ _00858_ _01539_ VPWR VGND _04678_ sg13g2_and2_1
X_10988_ _04678_ VPWR VGND _04679_ sg13g2_buf_1
X_10989_ _04674_ _04677_ _04679_ VPWR VGND _04680_ sg13g2_nand3_1
X_10990_ _00857_ _01536_ _01537_ VPWR VGND _04681_ sg13g2_nand3_1
X_10991_ _04681_ VPWR VGND _04682_ sg13g2_buf_1
X_10992_ _04674_ _04676_ _04682_ VPWR VGND _04683_ sg13g2_or3_1
X_10993_ _04667_ _04673_ _04680_ _04683_ VPWR VGND 
+ _04684_
+ sg13g2_a22oi_1
X_10994_ \atbs_core_0.dac_control_1.dac_counter_value[6]\ VPWR VGND _04685_ sg13g2_buf_1
X_10995_ _04685_ _04674_ _04677_ VPWR VGND _04686_ sg13g2_nand3_1
X_10996_ _04674_ _04685_ VPWR VGND _04687_ sg13g2_nor2b_1
X_10997_ _04677_ _04687_ VPWR VGND _04688_ sg13g2_nand2b_1
X_10998_ _04667_ _04673_ _04686_ _04688_ VPWR VGND 
+ _04689_
+ sg13g2_a22oi_1
X_10999_ _04685_ _04679_ VPWR VGND _04690_ sg13g2_nand2_1
X_11000_ \atbs_core_0.dac_control_1.dac_counter_value[5]\ VPWR VGND _04691_ sg13g2_buf_1
X_11001_ _04691_ _04677_ _04679_ VPWR VGND _04692_ sg13g2_nand3_1
X_11002_ _04685_ _04691_ _04677_ VPWR VGND _04693_ sg13g2_nand3_1
X_11003_ _04690_ _04692_ _04693_ VPWR VGND _04694_ sg13g2_nand3_1
X_11004_ _04626_ _04684_ _04689_ _04694_ VPWR VGND 
+ _04695_
+ sg13g2_nor4_2
X_11005_ _04622_ _01039_ _04625_ _04695_ VPWR VGND 
+ _04696_
+ sg13g2_nor4_1
X_11006_ \atbs_core_0.dac_control_1.dac_counter_value[8]\ _01039_ VPWR VGND _04697_ sg13g2_nor2_1
X_11007_ _04625_ _04695_ _04697_ VPWR VGND _04698_ sg13g2_o21ai_1
X_11008_ _00860_ _00858_ \atbs_core_0.adaptive_ctrl_0.spike_i\ VPWR VGND _04699_ sg13g2_a21oi_1
X_11009_ _01032_ _04699_ _00054_ VPWR VGND _04700_ sg13g2_a21oi_1
X_11010_ _04696_ _04698_ _04700_ VPWR VGND _04701_ sg13g2_nand3b_1
X_11011_ _04701_ VPWR VGND _04702_ sg13g2_buf_4
X_11012_ _04702_ VPWR VGND _04703_ sg13g2_buf_16
X_11013_ _04632_ _04649_ VPWR VGND _04704_ sg13g2_nand2_1
X_11014_ _01039_ _04699_ VPWR VGND _04705_ sg13g2_nor2_1
X_11015_ _04705_ VPWR VGND _04706_ sg13g2_buf_2
X_11016_ _04706_ VPWR VGND _04707_ sg13g2_buf_1
X_11017_ _00067_ VPWR VGND _04708_ sg13g2_buf_1
X_11018_ _04708_ _04649_ VPWR VGND _04709_ sg13g2_nand2_1
X_11019_ _04708_ _04649_ VPWR VGND _04710_ sg13g2_or2_1
X_11020_ _04709_ _04706_ _04710_ VPWR VGND _04711_ sg13g2_o21ai_1
X_11021_ _00068_ VPWR VGND _04712_ sg13g2_buf_1
X_11022_ _00858_ _01487_ VPWR VGND _04713_ sg13g2_nand2_1
X_11023_ _04708_ _00857_ _01453_ _01470_ VPWR VGND 
+ _04714_
+ sg13g2_nand4_1
X_11024_ _04708_ _00856_ VPWR VGND _04715_ sg13g2_nand2_1
X_11025_ _01231_ _01462_ _01450_ _01212_ _04715_ VPWR 
+ VGND
+ _04716_ sg13g2_a221oi_1
X_11026_ _01224_ _01498_ VPWR VGND _04717_ sg13g2_nand2_1
X_11027_ _04708_ _04382_ _04716_ _04717_ _04646_ VPWR 
+ VGND
+ _04718_ sg13g2_a221oi_1
X_11028_ _04357_ _04713_ _04714_ _04653_ _04718_ VPWR 
+ VGND
+ _04719_ sg13g2_a221oi_1
X_11029_ _00857_ _01487_ _04454_ VPWR VGND _04720_ sg13g2_a21oi_1
X_11030_ _00857_ _01487_ _04345_ _04355_ _00059_ VPWR 
+ VGND
+ _04721_ sg13g2_a221oi_1
X_11031_ _04720_ _04718_ _04721_ _04714_ _04651_ VPWR 
+ VGND
+ _04722_ sg13g2_a221oi_1
X_11032_ _00944_ _01462_ VPWR VGND _04723_ sg13g2_nor2_1
X_11033_ _00944_ _01498_ VPWR VGND _04724_ sg13g2_nor2_1
X_11034_ _01351_ _04723_ _04724_ _01344_ _04400_ VPWR 
+ VGND
+ _04725_ sg13g2_a221oi_1
X_11035_ _04725_ VPWR VGND _04726_ sg13g2_buf_1
X_11036_ _04669_ VPWR VGND _04727_ sg13g2_inv_1
X_11037_ _04658_ _04630_ _04726_ _04727_ VPWR VGND 
+ _04728_
+ sg13g2_a22oi_1
X_11038_ _04719_ _04722_ _04728_ VPWR VGND _04729_ sg13g2_o21ai_1
X_11039_ _04727_ _04726_ _04657_ VPWR VGND _04730_ sg13g2_a21oi_1
X_11040_ _04669_ _04664_ _04730_ VPWR VGND _04731_ sg13g2_a21oi_1
X_11041_ _04685_ _04682_ VPWR VGND _04732_ sg13g2_nand2_1
X_11042_ _04676_ _04732_ VPWR VGND _04733_ sg13g2_nand2_1
X_11043_ _04674_ _04732_ VPWR VGND _04734_ sg13g2_nand2_1
X_11044_ _04729_ _04731_ _04733_ _04734_ VPWR VGND 
+ _04735_
+ sg13g2_a22oi_1
X_11045_ _04674_ _04676_ _04732_ VPWR VGND _04736_ sg13g2_nand3_1
X_11046_ _04685_ _04682_ _04736_ VPWR VGND _04737_ sg13g2_o21ai_1
X_11047_ _04735_ _04737_ _04624_ VPWR VGND _04738_ sg13g2_o21ai_1
X_11048_ _04624_ _04735_ _04737_ VPWR VGND _04739_ sg13g2_nor3_1
X_11049_ _04623_ _04738_ _04739_ VPWR VGND _04740_ sg13g2_a21oi_2
X_11050_ _04712_ _04740_ VPWR VGND _04741_ sg13g2_nand2_1
X_11051_ _04704_ _04707_ _04711_ _04741_ VPWR VGND 
+ _04742_
+ sg13g2_a22oi_1
X_11052_ _04742_ _01036_ VPWR VGND _04743_ sg13g2_nand2b_1
X_11053_ _04632_ _04649_ VPWR VGND _04744_ sg13g2_nor2_1
X_11054_ _04632_ _04703_ VPWR VGND _04745_ sg13g2_nor2_2
X_11055_ _04703_ _04743_ _04744_ _04707_ _04745_ VPWR 
+ VGND
+ _00503_ sg13g2_a221oi_1
X_11056_ _04653_ _04646_ VPWR VGND _04746_ sg13g2_xnor2_1
X_11057_ _04709_ _04746_ VPWR VGND _04747_ sg13g2_xor2_1
X_11058_ _04712_ _04740_ _04706_ VPWR VGND _04748_ sg13g2_a21oi_2
X_11059_ _04647_ _04704_ VPWR VGND _04749_ sg13g2_xnor2_1
X_11060_ _04747_ _04748_ _04749_ _04707_ VPWR VGND 
+ _04750_
+ sg13g2_a22oi_1
X_11061_ _01037_ _04750_ VPWR VGND _04751_ sg13g2_nor2_1
X_11062_ \atbs_core_0.dac_control_1.dac_counter_value[1]\ _04751_ _04703_ VPWR VGND _00504_ sg13g2_mux2_1
X_11063_ _04632_ _04647_ _04649_ VPWR VGND _04752_ sg13g2_and3_1
X_11064_ _04654_ _04752_ VPWR VGND _04753_ sg13g2_or2_1
X_11065_ _04633_ _04753_ VPWR VGND _04754_ sg13g2_xnor2_1
X_11066_ _04653_ _04714_ _04718_ VPWR VGND _04755_ sg13g2_a21oi_1
X_11067_ _00058_ _04755_ VPWR VGND _04756_ sg13g2_xnor2_1
X_11068_ _04706_ _04756_ VPWR VGND _04757_ sg13g2_nor2_1
X_11069_ _04706_ _04754_ _04757_ _04741_ _04720_ VPWR 
+ VGND
+ _04758_ sg13g2_a221oi_1
X_11070_ _04633_ _04753_ VPWR VGND _04759_ sg13g2_xor2_1
X_11071_ _04707_ _04759_ _04748_ _04756_ _04652_ VPWR 
+ VGND
+ _04760_ sg13g2_a221oi_1
X_11072_ _01037_ _04758_ _04760_ VPWR VGND _04761_ sg13g2_nor3_1
X_11073_ _04633_ _04761_ _04703_ VPWR VGND _00505_ sg13g2_mux2_1
X_11074_ _04650_ _04655_ VPWR VGND _04762_ sg13g2_and2_1
X_11075_ _04657_ _04659_ VPWR VGND _04763_ sg13g2_and2_1
X_11076_ _04763_ VPWR VGND _04764_ sg13g2_buf_1
X_11077_ _04762_ _04764_ VPWR VGND _04765_ sg13g2_xor2_1
X_11078_ _04719_ _04722_ VPWR VGND _04766_ sg13g2_or2_1
X_11079_ _04764_ _04766_ VPWR VGND _04767_ sg13g2_xnor2_1
X_11080_ _04707_ _04765_ _04767_ _04748_ VPWR VGND 
+ _04768_
+ sg13g2_a22oi_1
X_11081_ _01037_ _04768_ VPWR VGND _04769_ sg13g2_nor2_1
X_11082_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ _04769_ _04703_ VPWR VGND _00506_ sg13g2_mux2_1
X_11083_ _04712_ _04740_ VPWR VGND _04770_ sg13g2_and2_1
X_11084_ _04770_ VPWR VGND _04771_ sg13g2_buf_2
X_11085_ _04658_ _04630_ VPWR VGND _04772_ sg13g2_nor2_1
X_11086_ _04659_ _04766_ _04772_ VPWR VGND _04773_ sg13g2_a21oi_1
X_11087_ _04727_ _04773_ VPWR VGND _04774_ sg13g2_xnor2_1
X_11088_ _04623_ _04624_ VPWR VGND _04775_ sg13g2_xor2_1
X_11089_ _04685_ _04682_ VPWR VGND _04776_ sg13g2_xor2_1
X_11090_ _04709_ _04710_ _04746_ _04776_ VPWR VGND 
+ _04777_
+ sg13g2_nand4_1
X_11091_ _00058_ _04720_ VPWR VGND _04778_ sg13g2_xnor2_1
X_11092_ _04712_ _04764_ _04778_ VPWR VGND _04779_ sg13g2_nand3_1
X_11093_ _04674_ _04676_ VPWR VGND _04780_ sg13g2_xor2_1
X_11094_ _04669_ _04726_ VPWR VGND _04781_ sg13g2_xnor2_1
X_11095_ _04780_ _04781_ VPWR VGND _04782_ sg13g2_nand2_1
X_11096_ _04775_ _04777_ _04779_ _04782_ VPWR VGND 
+ _04783_
+ sg13g2_nor4_1
X_11097_ _04706_ _04783_ VPWR VGND _04784_ sg13g2_or2_1
X_11098_ _04784_ VPWR VGND _04785_ sg13g2_buf_1
X_11099_ _04774_ _04785_ VPWR VGND _04786_ sg13g2_or2_1
X_11100_ _04631_ _04660_ VPWR VGND _04787_ sg13g2_nor2_1
X_11101_ _04662_ _04787_ VPWR VGND _04788_ sg13g2_xnor2_1
X_11102_ _04706_ _04788_ _04726_ VPWR VGND _04789_ sg13g2_a21oi_1
X_11103_ _04771_ _04786_ _04789_ VPWR VGND _04790_ sg13g2_o21ai_1
X_11104_ _04785_ _04774_ VPWR VGND _04791_ sg13g2_nand2b_1
X_11105_ _04661_ _04787_ VPWR VGND _04792_ sg13g2_xnor2_1
X_11106_ _04706_ _04792_ _04664_ VPWR VGND _04793_ sg13g2_a21oi_1
X_11107_ _04771_ _04791_ _04793_ VPWR VGND _04794_ sg13g2_o21ai_1
X_11108_ _01036_ _04702_ _04790_ _04794_ VPWR VGND 
+ _04795_
+ sg13g2_nand4_1
X_11109_ _04662_ _04703_ _04795_ VPWR VGND _00507_ sg13g2_o21ai_1
X_11110_ _04729_ _04731_ VPWR VGND _04796_ sg13g2_nand2_1
X_11111_ _04796_ _04780_ VPWR VGND _04797_ sg13g2_xnor2_1
X_11112_ _04667_ _04673_ VPWR VGND _04798_ sg13g2_nand2_1
X_11113_ _04798_ _04780_ VPWR VGND _04799_ sg13g2_xnor2_1
X_11114_ _04748_ _04797_ _04799_ _04707_ VPWR VGND 
+ _04800_
+ sg13g2_a22oi_1
X_11115_ _01037_ _04800_ VPWR VGND _04801_ sg13g2_nor2_1
X_11116_ _04691_ _04801_ _04703_ VPWR VGND _00508_ sg13g2_mux2_1
X_11117_ _04674_ _04677_ VPWR VGND _04802_ sg13g2_or2_1
X_11118_ _04674_ _04677_ VPWR VGND _04803_ sg13g2_nand2_1
X_11119_ _04667_ _04673_ _04802_ _04803_ VPWR VGND 
+ _04804_
+ sg13g2_a22oi_1
X_11120_ _04691_ _04677_ _04804_ VPWR VGND _04805_ sg13g2_a21oi_1
X_11121_ _04805_ _04776_ VPWR VGND _04806_ sg13g2_xnor2_1
X_11122_ _04806_ _04707_ VPWR VGND _04807_ sg13g2_nand2b_1
X_11123_ _04677_ _04796_ _04674_ VPWR VGND _04808_ sg13g2_a21o_1
X_11124_ _04677_ _04796_ _04808_ VPWR VGND _04809_ sg13g2_o21ai_1
X_11125_ _04809_ _04776_ VPWR VGND _04810_ sg13g2_xnor2_1
X_11126_ _04771_ _04706_ _04783_ _04810_ VPWR VGND 
+ _04811_
+ sg13g2_or4_1
X_11127_ _04807_ _04811_ _01037_ VPWR VGND _04812_ sg13g2_a21oi_1
X_11128_ _04685_ _04812_ _04703_ VPWR VGND _00509_ sg13g2_mux2_1
X_11129_ _04684_ _04689_ _04694_ VPWR VGND _04813_ sg13g2_nor3_1
X_11130_ _04813_ _04775_ VPWR VGND _04814_ sg13g2_xnor2_1
X_11131_ _04735_ _04737_ VPWR VGND _04815_ sg13g2_nor2_1
X_11132_ _04815_ _04775_ VPWR VGND _04816_ sg13g2_xor2_1
X_11133_ _04785_ _04816_ VPWR VGND _04817_ sg13g2_nor2_1
X_11134_ _04707_ _04814_ _04817_ _04741_ VPWR VGND 
+ _04818_
+ sg13g2_a22oi_1
X_11135_ \atbs_core_0.dac_control_1.dac_init_value[7]\ _01036_ VPWR VGND _04819_ sg13g2_nor2_1
X_11136_ _01036_ _04818_ _04819_ VPWR VGND _04820_ sg13g2_a21oi_1
X_11137_ _04623_ _04820_ _04703_ VPWR VGND _00510_ sg13g2_mux2_1
X_11138_ _04625_ _04695_ VPWR VGND _04821_ sg13g2_nor2_1
X_11139_ _04622_ _04821_ VPWR VGND _04822_ sg13g2_xnor2_1
X_11140_ _04712_ _04740_ _04707_ VPWR VGND _04823_ sg13g2_nor3_1
X_11141_ _04822_ _04707_ _04823_ VPWR VGND _04824_ sg13g2_a21oi_1
X_11142_ _01036_ _04703_ VPWR VGND _04825_ sg13g2_nand2_2
X_11143_ _04622_ _04702_ VPWR VGND _04826_ sg13g2_or2_1
X_11144_ _04824_ _04825_ _04826_ VPWR VGND _00511_ sg13g2_o21ai_1
X_11145_ \atbs_core_0.dac_control_1.dac_wr_o\ VPWR VGND _04827_ sg13g2_buf_1
X_11146_ dac_lower_o[0] _04632_ _04827_ VPWR VGND _00512_ sg13g2_mux2_1
X_11147_ dac_lower_o[1] \atbs_core_0.dac_control_1.dac_counter_value[1]\ _04827_ VPWR VGND _00513_ sg13g2_mux2_1
X_11148_ dac_lower_o[2] _04633_ _04827_ VPWR VGND _00514_ sg13g2_mux2_1
X_11149_ dac_lower_o[3] \atbs_core_0.dac_control_1.dac_counter_value[3]\ _04827_ VPWR VGND _00515_ sg13g2_mux2_1
X_11150_ dac_lower_o[4] _04661_ _04827_ VPWR VGND _00516_ sg13g2_mux2_1
X_11151_ dac_lower_o[5] _04691_ _04827_ VPWR VGND _00517_ sg13g2_mux2_1
X_11152_ dac_lower_o[6] _04685_ _04827_ VPWR VGND _00518_ sg13g2_mux2_1
X_11153_ dac_lower_o[7] _04623_ _04827_ VPWR VGND _00519_ sg13g2_mux2_1
X_11154_ \atbs_core_0.dac_control_1.n1727_q[1]\ \atbs_core_0.dac_control_1.n1727_q[0]\ VPWR VGND _04828_ sg13g2_nand2_1
X_11155_ _00053_ _04828_ VPWR VGND _04829_ sg13g2_or2_1
X_11156_ \atbs_core_0.dac_control_1.dac_change_in_progress\ _04829_ \atbs_core_0.dac_control_1.dac_counter_strb\ VPWR VGND _00520_ sg13g2_a21o_1
X_11157_ \atbs_core_0.debouncer_0.n1173_q[1]\ VPWR VGND _04830_ sg13g2_buf_1
X_11158_ \atbs_core_0.debouncer_0.n1173_q[0]\ VPWR VGND _04831_ sg13g2_buf_1
X_11159_ \atbs_core_0.debouncer_0.counter_value[1]\ VPWR VGND _04832_ sg13g2_buf_1
X_11160_ \atbs_core_0.debouncer_0.counter_value[0]\ VPWR VGND _04833_ sg13g2_buf_1
X_11161_ _04832_ _04833_ VPWR VGND _04834_ sg13g2_nor2b_1
X_11162_ \atbs_core_0.debouncer_0.counter_value[2]\ \atbs_core_0.debouncer_0.counter_value[3]\ _04834_ VPWR VGND _04835_ sg13g2_nand3b_1
X_11163_ _04835_ VPWR VGND _04836_ sg13g2_buf_1
X_11164_ \atbs_core_0.debouncer_0.bouncing_sync_d\ VPWR VGND _04837_ sg13g2_buf_1
X_11165_ _04837_ VPWR VGND _04838_ sg13g2_inv_1
X_11166_ _04831_ \atbs_core_0.debouncer_0.bouncing_sync\ _04838_ VPWR VGND _04839_ sg13g2_nor3_1
X_11167_ _04831_ _04836_ _04839_ VPWR VGND _04840_ sg13g2_a21oi_1
X_11168_ _04830_ _04840_ VPWR VGND _00521_ sg13g2_nor2_1
X_11169_ \atbs_core_0.debouncer_0.bouncing_sync\ VPWR VGND _04841_ sg13g2_inv_1
X_11170_ _04830_ _04841_ _04837_ VPWR VGND _04842_ sg13g2_nor3_1
X_11171_ _04830_ _04836_ _04842_ VPWR VGND _04843_ sg13g2_a21oi_1
X_11172_ _04831_ _04843_ VPWR VGND _00522_ sg13g2_nor2_1
X_11173_ _04831_ _04830_ VPWR VGND _04844_ sg13g2_xnor2_1
X_11174_ _04836_ _04844_ VPWR VGND _04845_ sg13g2_nor2_1
X_11175_ \atbs_core_0.debouncer_0.debounced\ _04837_ _04845_ VPWR VGND _00523_ sg13g2_mux2_1
X_11176_ \atbs_core_0.debouncer_1.n1173_q[1]\ VPWR VGND _04846_ sg13g2_buf_1
X_11177_ \atbs_core_0.debouncer_1.n1173_q[0]\ VPWR VGND _04847_ sg13g2_buf_1
X_11178_ \atbs_core_0.debouncer_1.counter_value[1]\ VPWR VGND _04848_ sg13g2_buf_1
X_11179_ \atbs_core_0.debouncer_1.counter_value[0]\ VPWR VGND _04849_ sg13g2_buf_1
X_11180_ _04848_ _04849_ VPWR VGND _04850_ sg13g2_nor2b_1
X_11181_ \atbs_core_0.debouncer_1.counter_value[2]\ \atbs_core_0.debouncer_1.counter_value[3]\ _04850_ VPWR VGND _04851_ sg13g2_nand3b_1
X_11182_ _04851_ VPWR VGND _04852_ sg13g2_buf_1
X_11183_ \atbs_core_0.debouncer_1.bouncing_sync_d\ VPWR VGND _04853_ sg13g2_buf_1
X_11184_ _04853_ VPWR VGND _04854_ sg13g2_inv_1
X_11185_ \atbs_core_0.debouncer_1.bouncing_sync\ _04854_ _04847_ VPWR VGND _04855_ sg13g2_nor3_1
X_11186_ _04847_ _04852_ _04855_ VPWR VGND _04856_ sg13g2_a21oi_1
X_11187_ _04846_ _04856_ VPWR VGND _00524_ sg13g2_nor2_1
X_11188_ \atbs_core_0.debouncer_1.bouncing_sync\ VPWR VGND _04857_ sg13g2_inv_1
X_11189_ _04857_ _04853_ _04846_ VPWR VGND _04858_ sg13g2_nor3_1
X_11190_ _04846_ _04852_ _04858_ VPWR VGND _04859_ sg13g2_a21oi_1
X_11191_ _04847_ _04859_ VPWR VGND _00525_ sg13g2_nor2_1
X_11192_ _04847_ _04846_ VPWR VGND _04860_ sg13g2_xnor2_1
X_11193_ _04852_ _04860_ VPWR VGND _04861_ sg13g2_nor2_1
X_11194_ \atbs_core_0.adaptive_mode_debounced\ _04853_ _04861_ VPWR VGND _00526_ sg13g2_mux2_1
X_11195_ \atbs_core_0.debouncer_2.n1173_q[1]\ VPWR VGND _04862_ sg13g2_buf_1
X_11196_ \atbs_core_0.debouncer_2.n1173_q[0]\ VPWR VGND _04863_ sg13g2_buf_1
X_11197_ \atbs_core_0.debouncer_2.counter_value[1]\ VPWR VGND _04864_ sg13g2_buf_1
X_11198_ \atbs_core_0.debouncer_2.counter_value[0]\ VPWR VGND _04865_ sg13g2_buf_1
X_11199_ _04864_ _04865_ VPWR VGND _04866_ sg13g2_nor2b_1
X_11200_ \atbs_core_0.debouncer_2.counter_value[2]\ \atbs_core_0.debouncer_2.counter_value[3]\ _04866_ VPWR VGND _04867_ sg13g2_nand3b_1
X_11201_ _04867_ VPWR VGND _04868_ sg13g2_buf_1
X_11202_ \atbs_core_0.debouncer_2.bouncing_sync_d\ VPWR VGND _04869_ sg13g2_buf_1
X_11203_ _04869_ VPWR VGND _04870_ sg13g2_inv_1
X_11204_ \atbs_core_0.debouncer_2.bouncing_sync\ _04870_ _04863_ VPWR VGND _04871_ sg13g2_nor3_1
X_11205_ _04863_ _04868_ _04871_ VPWR VGND _04872_ sg13g2_a21oi_1
X_11206_ _04862_ _04872_ VPWR VGND _00527_ sg13g2_nor2_1
X_11207_ \atbs_core_0.debouncer_2.bouncing_sync\ VPWR VGND _04873_ sg13g2_inv_1
X_11208_ _04873_ _04869_ _04862_ VPWR VGND _04874_ sg13g2_nor3_1
X_11209_ _04862_ _04868_ _04874_ VPWR VGND _04875_ sg13g2_a21oi_1
X_11210_ _04863_ _04875_ VPWR VGND _00528_ sg13g2_nor2_1
X_11211_ _04863_ _04862_ VPWR VGND _04876_ sg13g2_xnor2_1
X_11212_ _04868_ _04876_ VPWR VGND _04877_ sg13g2_nor2_1
X_11213_ _00853_ _04869_ _04877_ VPWR VGND _00529_ sg13g2_mux2_1
X_11214_ \atbs_core_0.debouncer_3.n1173_q[1]\ VPWR VGND _04878_ sg13g2_buf_1
X_11215_ \atbs_core_0.debouncer_3.n1173_q[0]\ VPWR VGND _04879_ sg13g2_buf_1
X_11216_ \atbs_core_0.debouncer_3.counter_value[1]\ VPWR VGND _04880_ sg13g2_buf_1
X_11217_ \atbs_core_0.debouncer_3.counter_value[0]\ VPWR VGND _04881_ sg13g2_buf_1
X_11218_ _04880_ _04881_ VPWR VGND _04882_ sg13g2_nor2b_1
X_11219_ \atbs_core_0.debouncer_3.counter_value[2]\ \atbs_core_0.debouncer_3.counter_value[3]\ _04882_ VPWR VGND _04883_ sg13g2_nand3b_1
X_11220_ _04883_ VPWR VGND _04884_ sg13g2_buf_1
X_11221_ \atbs_core_0.debouncer_3.bouncing_sync_d\ VPWR VGND _04885_ sg13g2_buf_1
X_11222_ _04885_ VPWR VGND _04886_ sg13g2_inv_1
X_11223_ \atbs_core_0.debouncer_3.bouncing_sync\ _04886_ _04879_ VPWR VGND _04887_ sg13g2_nor3_1
X_11224_ _04879_ _04884_ _04887_ VPWR VGND _04888_ sg13g2_a21oi_1
X_11225_ _04878_ _04888_ VPWR VGND _00530_ sg13g2_nor2_1
X_11226_ \atbs_core_0.debouncer_3.bouncing_sync\ VPWR VGND _04889_ sg13g2_inv_1
X_11227_ _04889_ _04885_ _04878_ VPWR VGND _04890_ sg13g2_nor3_1
X_11228_ _04878_ _04884_ _04890_ VPWR VGND _04891_ sg13g2_a21oi_1
X_11229_ _04879_ _04891_ VPWR VGND _00531_ sg13g2_nor2_1
X_11230_ _04878_ _04879_ VPWR VGND _04892_ sg13g2_xnor2_1
X_11231_ _04884_ _04892_ VPWR VGND _04893_ sg13g2_nor2_1
X_11232_ \atbs_core_0.debouncer_3.debounced\ _04885_ _04893_ VPWR VGND _00532_ sg13g2_mux2_1
X_11233_ \atbs_core_0.debouncer_4.n1173_q[1]\ VPWR VGND _04894_ sg13g2_buf_1
X_11234_ \atbs_core_0.debouncer_4.n1173_q[0]\ VPWR VGND _04895_ sg13g2_buf_1
X_11235_ \atbs_core_0.debouncer_4.counter_value[1]\ VPWR VGND _04896_ sg13g2_buf_1
X_11236_ \atbs_core_0.debouncer_4.counter_value[0]\ VPWR VGND _04897_ sg13g2_buf_1
X_11237_ _04896_ _04897_ VPWR VGND _04898_ sg13g2_nor2b_1
X_11238_ \atbs_core_0.debouncer_4.counter_value[2]\ \atbs_core_0.debouncer_4.counter_value[3]\ _04898_ VPWR VGND _04899_ sg13g2_nand3b_1
X_11239_ _04899_ VPWR VGND _04900_ sg13g2_buf_1
X_11240_ \atbs_core_0.debouncer_4.bouncing_sync_d\ VPWR VGND _04901_ sg13g2_buf_1
X_11241_ _04901_ VPWR VGND _04902_ sg13g2_inv_1
X_11242_ \atbs_core_0.debouncer_4.bouncing_sync\ _04902_ _04895_ VPWR VGND _04903_ sg13g2_nor3_1
X_11243_ _04895_ _04900_ _04903_ VPWR VGND _04904_ sg13g2_a21oi_1
X_11244_ _04894_ _04904_ VPWR VGND _00533_ sg13g2_nor2_1
X_11245_ \atbs_core_0.debouncer_4.bouncing_sync\ VPWR VGND _04905_ sg13g2_inv_1
X_11246_ _04905_ _04901_ _04894_ VPWR VGND _04906_ sg13g2_nor3_1
X_11247_ _04894_ _04900_ _04906_ VPWR VGND _04907_ sg13g2_a21oi_1
X_11248_ _04895_ _04907_ VPWR VGND _00534_ sg13g2_nor2_1
X_11249_ _04895_ _04894_ VPWR VGND _04908_ sg13g2_xnor2_1
X_11250_ _04900_ _04908_ VPWR VGND _04909_ sg13g2_nor2_1
X_11251_ \atbs_core_0.debouncer_4.debounced\ _04901_ _04909_ VPWR VGND _00535_ sg13g2_mux2_1
X_11252_ \atbs_core_0.debouncer_5.n1173_q[1]\ VPWR VGND _04910_ sg13g2_buf_1
X_11253_ \atbs_core_0.debouncer_5.n1173_q[0]\ VPWR VGND _04911_ sg13g2_buf_1
X_11254_ \atbs_core_0.debouncer_5.counter_value[1]\ VPWR VGND _04912_ sg13g2_buf_1
X_11255_ \atbs_core_0.debouncer_5.counter_value[0]\ VPWR VGND _04913_ sg13g2_buf_1
X_11256_ _04912_ _04913_ VPWR VGND _04914_ sg13g2_nor2b_1
X_11257_ \atbs_core_0.debouncer_5.counter_value[2]\ \atbs_core_0.debouncer_5.counter_value[3]\ _04914_ VPWR VGND _04915_ sg13g2_nand3b_1
X_11258_ _04915_ VPWR VGND _04916_ sg13g2_buf_1
X_11259_ \atbs_core_0.debouncer_5.bouncing_sync_d\ VPWR VGND _04917_ sg13g2_buf_1
X_11260_ _04917_ VPWR VGND _04918_ sg13g2_inv_1
X_11261_ _04911_ \atbs_core_0.debouncer_5.bouncing_sync\ _04918_ VPWR VGND _04919_ sg13g2_nor3_1
X_11262_ _04911_ _04916_ _04919_ VPWR VGND _04920_ sg13g2_a21oi_1
X_11263_ _04910_ _04920_ VPWR VGND _00536_ sg13g2_nor2_1
X_11264_ \atbs_core_0.debouncer_5.bouncing_sync\ VPWR VGND _04921_ sg13g2_inv_1
X_11265_ _04910_ _04921_ _04917_ VPWR VGND _04922_ sg13g2_nor3_1
X_11266_ _04910_ _04916_ _04922_ VPWR VGND _04923_ sg13g2_a21oi_1
X_11267_ _04911_ _04923_ VPWR VGND _00537_ sg13g2_nor2_1
X_11268_ _04911_ _04910_ VPWR VGND _04924_ sg13g2_xnor2_1
X_11269_ _04916_ _04924_ VPWR VGND _04925_ sg13g2_nor2_1
X_11270_ \atbs_core_0.debouncer_5.debounced\ _04917_ _04925_ VPWR VGND _00538_ sg13g2_mux2_1
X_11271_ \atbs_core_0.memory2uart_0.tx_strb_i\ VPWR VGND _04926_ sg13g2_inv_1
X_11272_ \atbs_core_0.memory2uart_0.read_strb_i\ VPWR VGND _04927_ sg13g2_buf_1
X_11273_ _04927_ VPWR VGND _04928_ sg13g2_inv_1
X_11274_ _04926_ \atbs_core_0.memory2uart_0.counter[1]\ _04928_ VPWR VGND \atbs_core_0.memory2uart_0.n2023_o\ sg13g2_o21ai_1
X_11275_ _04927_ VPWR VGND _04929_ sg13g2_buf_1
X_11276_ _04929_ VPWR VGND _04930_ sg13g2_buf_1
X_11277_ _04926_ \atbs_core_0.memory2uart_0.counter[1]\ VPWR VGND _04931_ sg13g2_nor2_1
X_11278_ _04931_ VPWR VGND _04932_ sg13g2_buf_1
X_11279_ _04932_ VPWR VGND _04933_ sg13g2_buf_1
X_11280_ _04932_ VPWR VGND _04934_ sg13g2_buf_1
X_11281_ _04934_ \atbs_core_0.uart_0.uart_tx_0.n2783_o\ VPWR VGND _04935_ sg13g2_nor2b_1
X_11282_ \atbs_core_0.memory2uart_0.n2009_o[0]\ _04933_ _04935_ VPWR VGND _04936_ sg13g2_a21oi_1
X_11283_ _04929_ VPWR VGND _04937_ sg13g2_buf_1
X_11284_ _04937_ \atbs_core_0.b_data[16]\ VPWR VGND _04938_ sg13g2_nand2_1
X_11285_ _04930_ _04936_ _04938_ VPWR VGND _00539_ sg13g2_o21ai_1
X_11286_ _04934_ \atbs_core_0.memory2uart_0.n2009_o[2]\ VPWR VGND _04939_ sg13g2_nor2b_1
X_11287_ \atbs_core_0.memory2uart_0.n2009_o[10]\ _04933_ _04939_ VPWR VGND _04940_ sg13g2_a21oi_1
X_11288_ _04937_ \atbs_core_0.b_data[10]\ VPWR VGND _04941_ sg13g2_nand2_1
X_11289_ _04930_ _04940_ _04941_ VPWR VGND _00540_ sg13g2_o21ai_1
X_11290_ _04932_ VPWR VGND _04942_ sg13g2_buf_1
X_11291_ _04934_ \atbs_core_0.memory2uart_0.n2009_o[3]\ VPWR VGND _04943_ sg13g2_nor2b_1
X_11292_ \atbs_core_0.memory2uart_0.n2009_o[11]\ _04942_ _04943_ VPWR VGND _04944_ sg13g2_a21oi_1
X_11293_ _04929_ \atbs_core_0.b_data[11]\ VPWR VGND _04945_ sg13g2_nand2_1
X_11294_ _04930_ _04944_ _04945_ VPWR VGND _00541_ sg13g2_o21ai_1
X_11295_ _04934_ \atbs_core_0.memory2uart_0.n2009_o[4]\ VPWR VGND _04946_ sg13g2_nor2b_1
X_11296_ \atbs_core_0.memory2uart_0.n2009_o[12]\ _04942_ _04946_ VPWR VGND _04947_ sg13g2_a21oi_1
X_11297_ _04929_ \atbs_core_0.b_data[12]\ VPWR VGND _04948_ sg13g2_nand2_1
X_11298_ _04930_ _04947_ _04948_ VPWR VGND _00542_ sg13g2_o21ai_1
X_11299_ _04934_ \atbs_core_0.memory2uart_0.n2009_o[5]\ VPWR VGND _04949_ sg13g2_nor2b_1
X_11300_ \atbs_core_0.memory2uart_0.n2009_o[13]\ _04942_ _04949_ VPWR VGND _04950_ sg13g2_a21oi_1
X_11301_ _04929_ \atbs_core_0.b_data[13]\ VPWR VGND _04951_ sg13g2_nand2_1
X_11302_ _04930_ _04950_ _04951_ VPWR VGND _00543_ sg13g2_o21ai_1
X_11303_ _04934_ \atbs_core_0.memory2uart_0.n2009_o[6]\ VPWR VGND _04952_ sg13g2_nor2b_1
X_11304_ \atbs_core_0.memory2uart_0.n2009_o[14]\ _04942_ _04952_ VPWR VGND _04953_ sg13g2_a21oi_1
X_11305_ _04929_ \atbs_core_0.b_data[14]\ VPWR VGND _04954_ sg13g2_nand2_1
X_11306_ _04930_ _04953_ _04954_ VPWR VGND _00544_ sg13g2_o21ai_1
X_11307_ _04932_ \atbs_core_0.memory2uart_0.n2009_o[7]\ VPWR VGND _04955_ sg13g2_nor2b_1
X_11308_ \atbs_core_0.memory2uart_0.n2009_o[15]\ _04942_ _04955_ VPWR VGND _04956_ sg13g2_a21oi_1
X_11309_ _04929_ \atbs_core_0.b_data[15]\ VPWR VGND _04957_ sg13g2_nand2_1
X_11310_ _04930_ _04956_ _04957_ VPWR VGND _00545_ sg13g2_o21ai_1
X_11311_ \atbs_core_0.memory2uart_0.n2009_o[8]\ \atbs_core_0.b_data[0]\ _04937_ VPWR VGND _00546_ sg13g2_mux2_1
X_11312_ \atbs_core_0.memory2uart_0.n2009_o[9]\ \atbs_core_0.b_data[1]\ _04937_ VPWR VGND _00547_ sg13g2_mux2_1
X_11313_ \atbs_core_0.memory2uart_0.n2009_o[10]\ \atbs_core_0.b_data[2]\ _04937_ VPWR VGND _00548_ sg13g2_mux2_1
X_11314_ \atbs_core_0.memory2uart_0.n2009_o[11]\ \atbs_core_0.b_data[3]\ _04937_ VPWR VGND _00549_ sg13g2_mux2_1
X_11315_ _04932_ \atbs_core_0.uart_0.uart_tx_0.n2784_o\ VPWR VGND _04958_ sg13g2_nor2b_1
X_11316_ \atbs_core_0.memory2uart_0.n2009_o[1]\ _04942_ _04958_ VPWR VGND _04959_ sg13g2_a21oi_1
X_11317_ _04929_ \atbs_core_0.b_data[17]\ VPWR VGND _04960_ sg13g2_nand2_1
X_11318_ _04930_ _04959_ _04960_ VPWR VGND _00550_ sg13g2_o21ai_1
X_11319_ \atbs_core_0.memory2uart_0.n2009_o[12]\ \atbs_core_0.b_data[4]\ _04937_ VPWR VGND _00551_ sg13g2_mux2_1
X_11320_ \atbs_core_0.memory2uart_0.n2009_o[13]\ \atbs_core_0.b_data[5]\ _04937_ VPWR VGND _00552_ sg13g2_mux2_1
X_11321_ \atbs_core_0.memory2uart_0.n2009_o[14]\ \atbs_core_0.b_data[6]\ _04937_ VPWR VGND _00553_ sg13g2_mux2_1
X_11322_ \atbs_core_0.memory2uart_0.n2009_o[15]\ \atbs_core_0.b_data[7]\ _04937_ VPWR VGND _00554_ sg13g2_mux2_1
X_11323_ \atbs_core_0.memory2uart_0.n2009_o[2]\ _04942_ VPWR VGND _04961_ sg13g2_nand2b_1
X_11324_ \atbs_core_0.uart_0.uart_tx_0.n2785_o\ _04933_ _04961_ VPWR VGND _04962_ sg13g2_o21ai_1
X_11325_ _04928_ \atbs_core_0.b_data[18]\ VPWR VGND _04963_ sg13g2_nor2_1
X_11326_ _04928_ _04962_ _04963_ VPWR VGND _00555_ sg13g2_a21oi_1
X_11327_ \atbs_core_0.memory2uart_0.n2009_o[3]\ _04942_ VPWR VGND _04964_ sg13g2_nand2b_1
X_11328_ \atbs_core_0.uart_0.uart_tx_0.n2786_o\ _04933_ _04964_ VPWR VGND _04965_ sg13g2_o21ai_1
X_11329_ _04928_ _04965_ _04963_ VPWR VGND _00556_ sg13g2_a21oi_1
X_11330_ \atbs_core_0.memory2uart_0.n2009_o[4]\ _04934_ VPWR VGND _04966_ sg13g2_nand2b_1
X_11331_ \atbs_core_0.uart_0.uart_tx_0.n2787_o\ _04933_ _04966_ VPWR VGND _04967_ sg13g2_o21ai_1
X_11332_ _04928_ _04967_ _04963_ VPWR VGND _00557_ sg13g2_a21oi_1
X_11333_ \atbs_core_0.memory2uart_0.n2009_o[5]\ _04934_ VPWR VGND _04968_ sg13g2_nand2b_1
X_11334_ \atbs_core_0.uart_0.uart_tx_0.n2788_o\ _04933_ _04968_ VPWR VGND _04969_ sg13g2_o21ai_1
X_11335_ _04928_ _04969_ _04963_ VPWR VGND _00558_ sg13g2_a21oi_1
X_11336_ \atbs_core_0.memory2uart_0.n2009_o[6]\ _04934_ VPWR VGND _04970_ sg13g2_nand2b_1
X_11337_ \atbs_core_0.uart_0.uart_tx_0.n2789_o\ _04933_ _04970_ VPWR VGND _04971_ sg13g2_o21ai_1
X_11338_ _04928_ _04971_ _04963_ VPWR VGND _00559_ sg13g2_a21oi_1
X_11339_ \atbs_core_0.memory2uart_0.n2009_o[7]\ _04934_ VPWR VGND _04972_ sg13g2_nand2b_1
X_11340_ \atbs_core_0.uart_0.uart_tx_0.n2790_o\ _04933_ _04972_ VPWR VGND _04973_ sg13g2_o21ai_1
X_11341_ _04928_ _04973_ _04963_ VPWR VGND _00560_ sg13g2_a21oi_1
X_11342_ _04932_ \atbs_core_0.memory2uart_0.n2009_o[0]\ VPWR VGND _04974_ sg13g2_nor2b_1
X_11343_ \atbs_core_0.memory2uart_0.n2009_o[8]\ _04942_ _04974_ VPWR VGND _04975_ sg13g2_a21oi_1
X_11344_ _04929_ \atbs_core_0.b_data[8]\ VPWR VGND _04976_ sg13g2_nand2_1
X_11345_ _04930_ _04975_ _04976_ VPWR VGND _00561_ sg13g2_o21ai_1
X_11346_ _04932_ \atbs_core_0.memory2uart_0.n2009_o[1]\ VPWR VGND _04977_ sg13g2_nor2b_1
X_11347_ \atbs_core_0.memory2uart_0.n2009_o[9]\ _04942_ _04977_ VPWR VGND _04978_ sg13g2_a21oi_1
X_11348_ _04929_ \atbs_core_0.b_data[9]\ VPWR VGND _04979_ sg13g2_nand2_1
X_11349_ _04930_ _04978_ _04979_ VPWR VGND _00562_ sg13g2_o21ai_1
X_11350_ _04933_ _04926_ \atbs_core_0.memory2uart_0.counter[0]\ VPWR VGND _00563_ sg13g2_mux2_1
X_11351_ \atbs_core_0.memory2uart_0.tx_strb_i\ \atbs_core_0.memory2uart_0.counter[1]\ VPWR VGND _04980_ sg13g2_nor2b_1
X_11352_ \atbs_core_0.memory2uart_0.counter[0]\ _04933_ _04980_ VPWR VGND _00564_ sg13g2_a21o_1
X_11353_ \atbs_core_0.detection_en\ VPWR VGND _04981_ sg13g2_inv_1
X_11354_ _01069_ _00842_ VPWR VGND _04982_ sg13g2_nor2_1
X_11355_ _04981_ _04982_ _01185_ VPWR VGND _00565_ sg13g2_o21ai_1
X_11356_ _00986_ _00984_ VPWR VGND _04983_ sg13g2_nor2_1
X_11357_ _00984_ _00987_ _04983_ _00985_ VPWR VGND 
+ _04984_
+ sg13g2_a22oi_1
X_11358_ _00842_ VPWR VGND _04985_ sg13g2_buf_1
X_11359_ _01069_ _04985_ _00843_ VPWR VGND _04986_ sg13g2_nand3_1
X_11360_ _04984_ _04986_ VPWR VGND _04987_ sg13g2_nor2_1
X_11361_ _04985_ \atbs_core_0.n1056_q\ _01069_ VPWR VGND _04988_ sg13g2_a21oi_1
X_11362_ _00844_ _01092_ VPWR VGND _04989_ sg13g2_nand2_1
X_11363_ _04985_ _04989_ \atbs_core_0.n1056_q\ VPWR VGND _04990_ sg13g2_a21oi_1
X_11364_ _04987_ _04988_ _04990_ VPWR VGND _00566_ sg13g2_nor3_1
X_11365_ _00989_ _04986_ VPWR VGND _04991_ sg13g2_or2_1
X_11366_ _00845_ _04982_ VPWR VGND _04992_ sg13g2_nand2_1
X_11367_ _00982_ _04991_ _04992_ _00989_ VPWR VGND 
+ _00567_
+ sg13g2_a22oi_1
X_11368_ \atbs_core_0.analog_trigger_uart\ VPWR VGND _04993_ sg13g2_inv_1
X_11369_ _01046_ VPWR VGND _04994_ sg13g2_inv_1
X_11370_ _01042_ \atbs_core_0.n1061_q\ VPWR VGND _04995_ sg13g2_nor2_1
X_11371_ _00050_ _04995_ VPWR VGND _04996_ sg13g2_nand2_1
X_11372_ _01077_ \atbs_core_0.n1067_q\ VPWR VGND _04997_ sg13g2_or2_1
X_11373_ _04994_ _04996_ _04997_ VPWR VGND _04998_ sg13g2_nor3_1
X_11374_ _01087_ _01055_ VPWR VGND _04999_ sg13g2_and2_1
X_11375_ _04999_ VPWR VGND _05000_ sg13g2_buf_1
X_11376_ _01050_ _04998_ _05000_ VPWR VGND _05001_ sg13g2_nand3_1
X_11377_ \atbs_core_0.uart_0.rx_data_strb_o\ _04993_ _05001_ VPWR VGND _00568_ sg13g2_o21ai_1
X_11378_ _01051_ _01053_ _01052_ VPWR VGND _05002_ sg13g2_o21ai_1
X_11379_ _01058_ _05002_ VPWR VGND _05003_ sg13g2_nand2b_1
X_11380_ _01050_ _05003_ VPWR VGND _05004_ sg13g2_and2_1
X_11381_ \atbs_core_0.uart_0.uart_rx_0.n2917_o\ \atbs_core_0.uart_0.uart_rx_0.n2915_o\ _01045_ VPWR VGND _05005_ sg13g2_nor3_1
X_11382_ _01076_ _00048_ _05004_ _05005_ VPWR VGND 
+ _05006_
+ sg13g2_nand4_1
X_11383_ _01043_ _01088_ VPWR VGND _05007_ sg13g2_nand2_1
X_11384_ _01042_ \atbs_core_0.analog_trigger_uart\ \atbs_core_0.n1061_q\ VPWR VGND _05008_ sg13g2_o21ai_1
X_11385_ _05006_ _05007_ _05008_ VPWR VGND _00569_ sg13g2_o21ai_1
X_11386_ _01048_ _01083_ _04996_ _05006_ VPWR VGND 
+ _05009_
+ sg13g2_nor4_1
X_11387_ _01077_ _04996_ _05009_ VPWR VGND _00570_ sg13g2_a21o_1
X_11388_ _01056_ \atbs_core_0.uart_0.uart_rx_0.n2915_o\ _01045_ VPWR VGND _05010_ sg13g2_nor3_1
X_11389_ _05010_ VPWR VGND _05011_ sg13g2_buf_1
X_11390_ _01084_ _05011_ VPWR VGND _05012_ sg13g2_and2_1
X_11391_ _05012_ VPWR VGND _05013_ sg13g2_buf_1
X_11392_ _01048_ _01082_ _05011_ VPWR VGND _05014_ sg13g2_nand3_1
X_11393_ _05014_ VPWR VGND _05015_ sg13g2_buf_1
X_11394_ _05013_ _05015_ VPWR VGND _05016_ sg13g2_nand2b_1
X_11395_ _05000_ _05011_ VPWR VGND _05017_ sg13g2_nand2_1
X_11396_ _05016_ _05017_ VPWR VGND _05018_ sg13g2_nand2b_1
X_11397_ _05018_ VPWR VGND _05019_ sg13g2_buf_1
X_11398_ _01077_ _00050_ _04995_ _05019_ VPWR VGND 
+ _05020_
+ sg13g2_nand4_1
X_11399_ _05020_ VPWR VGND _05021_ sg13g2_buf_1
X_11400_ _05013_ _00105_ _05021_ VPWR VGND _00571_ sg13g2_mux2_1
X_11401_ _00106_ VPWR VGND _05022_ sg13g2_inv_1
X_11402_ _05016_ _05021_ VPWR VGND _05023_ sg13g2_nor2_1
X_11403_ _05022_ _05021_ _05023_ VPWR VGND _00572_ sg13g2_a21oi_1
X_11404_ _01088_ _05011_ VPWR VGND _05024_ sg13g2_and2_1
X_11405_ _05024_ VPWR VGND _05025_ sg13g2_buf_1
X_11406_ _05025_ _00767_ _05021_ VPWR VGND _00573_ sg13g2_mux2_1
X_11407_ _05013_ _00762_ _05021_ VPWR VGND _00574_ sg13g2_mux2_1
X_11408_ _01051_ _05015_ VPWR VGND _05026_ sg13g2_nor2_1
X_11409_ _05026_ _00754_ _05021_ VPWR VGND _00575_ sg13g2_mux2_1
X_11410_ _00107_ _05021_ VPWR VGND _05027_ sg13g2_nand2_1
X_11411_ _05015_ _05021_ _05027_ VPWR VGND _00576_ sg13g2_o21ai_1
X_11412_ _00780_ _05021_ _05023_ VPWR VGND _00577_ sg13g2_a21oi_1
X_11413_ _00049_ _01046_ VPWR VGND _05028_ sg13g2_and2_1
X_11414_ _01051_ _01054_ VPWR VGND _05029_ sg13g2_and2_1
X_11415_ _05029_ VPWR VGND _05030_ sg13g2_buf_1
X_11416_ _01087_ _05030_ VPWR VGND _05031_ sg13g2_and2_1
X_11417_ _01078_ _05028_ _05004_ _05031_ VPWR VGND 
+ _05032_
+ sg13g2_nand4_1
X_11418_ _01076_ _01078_ _05032_ VPWR VGND _00578_ sg13g2_o21ai_1
X_11419_ _01048_ _01055_ _05011_ VPWR VGND _05033_ sg13g2_and3_1
X_11420_ _05033_ VPWR VGND _05034_ sg13g2_buf_1
X_11421_ \atbs_core_0.n1067_q\ _01078_ VPWR VGND _05035_ sg13g2_and2_1
X_11422_ _05035_ VPWR VGND _05036_ sg13g2_buf_1
X_11423_ _05019_ _05034_ _05036_ VPWR VGND _05037_ sg13g2_o21ai_1
X_11424_ _05037_ VPWR VGND _05038_ sg13g2_buf_1
X_11425_ _05026_ \atbs_core_0.n1068_q[1]\ _05038_ VPWR VGND _00579_ sg13g2_mux2_1
X_11426_ _05013_ _04355_ _05038_ VPWR VGND _00580_ sg13g2_mux2_1
X_11427_ _00108_ _05038_ VPWR VGND _05039_ sg13g2_nand2_1
X_11428_ _05025_ _05038_ _05039_ VPWR VGND _00581_ sg13g2_o21ai_1
X_11429_ \atbs_core_0.n1068_q[4]\ _05038_ VPWR VGND _05040_ sg13g2_nand2_1
X_11430_ _05017_ _05038_ _05040_ VPWR VGND _00582_ sg13g2_o21ai_1
X_11431_ _05034_ _05036_ \atbs_core_0.n1068_q[5]\ VPWR VGND _05041_ sg13g2_a21oi_1
X_11432_ _05019_ _05036_ _05041_ VPWR VGND _00583_ sg13g2_a21oi_1
X_11433_ _01048_ _00077_ _04998_ _05030_ VPWR VGND 
+ _05042_
+ sg13g2_nand4_1
X_11434_ _04996_ _04997_ _01049_ VPWR VGND _05043_ sg13g2_o21ai_1
X_11435_ _01049_ _05042_ _05043_ VPWR VGND _00584_ sg13g2_o21ai_1
X_11436_ _05016_ _05034_ VPWR VGND _05044_ sg13g2_nor2_1
X_11437_ _05019_ _05034_ VPWR VGND _05045_ sg13g2_nor2_1
X_11438_ _05011_ _05031_ VPWR VGND _05046_ sg13g2_nand2_1
X_11439_ _01049_ _01080_ VPWR VGND _05047_ sg13g2_nand2_1
X_11440_ _05045_ _05046_ _05047_ VPWR VGND _05048_ sg13g2_a21oi_1
X_11441_ _05048_ VPWR VGND _05049_ sg13g2_buf_1
X_11442_ _05049_ VPWR VGND _05050_ sg13g2_buf_1
X_11443_ _00109_ _05044_ _05050_ VPWR VGND _00585_ sg13g2_mux2_1
X_11444_ _00110_ _05034_ _05049_ VPWR VGND _00586_ sg13g2_mux2_1
X_11445_ _00111_ VPWR VGND _05051_ sg13g2_inv_1
X_11446_ _05045_ _05049_ VPWR VGND _05052_ sg13g2_nand2_1
X_11447_ _05051_ _05050_ _05052_ VPWR VGND _00587_ sg13g2_o21ai_1
X_11448_ _00112_ VPWR VGND _05053_ sg13g2_inv_1
X_11449_ _05026_ _05049_ VPWR VGND _05054_ sg13g2_nand2_1
X_11450_ _05053_ _05050_ _05054_ VPWR VGND _00588_ sg13g2_o21ai_1
X_11451_ _05013_ _05026_ VPWR VGND _05055_ sg13g2_nor2_1
X_11452_ _00113_ _05049_ VPWR VGND _05056_ sg13g2_nor2_1
X_11453_ _05050_ _05055_ _05056_ VPWR VGND _00589_ sg13g2_a21oi_1
X_11454_ _05016_ _05049_ VPWR VGND _05057_ sg13g2_nand2b_1
X_11455_ _01674_ _05050_ _05057_ VPWR VGND _00590_ sg13g2_o21ai_1
X_11456_ _05019_ _05049_ VPWR VGND _05058_ sg13g2_nand2b_1
X_11457_ _02491_ _05050_ _05058_ VPWR VGND _00591_ sg13g2_o21ai_1
X_11458_ _01697_ _05050_ _05052_ VPWR VGND _00592_ sg13g2_o21ai_1
X_11459_ _03714_ _05050_ _05054_ VPWR VGND _00593_ sg13g2_o21ai_1
X_11460_ _05013_ _05049_ VPWR VGND _05059_ sg13g2_nand2_1
X_11461_ _01780_ _05050_ _05059_ VPWR VGND _00594_ sg13g2_o21ai_1
X_11462_ _00114_ _05015_ _05049_ VPWR VGND _00595_ sg13g2_mux2_1
X_11463_ _05017_ _05055_ VPWR VGND _05060_ sg13g2_nand2_1
X_11464_ _05049_ _05060_ VPWR VGND _05061_ sg13g2_nand2_1
X_11465_ _01744_ _05050_ _05061_ VPWR VGND _00596_ sg13g2_o21ai_1
X_11466_ _00077_ _01081_ _05000_ _05005_ VPWR VGND 
+ _05062_
+ sg13g2_nand4_1
X_11467_ _01075_ _01081_ _05062_ VPWR VGND _00597_ sg13g2_o21ai_1
X_11468_ _01081_ VPWR VGND _05063_ sg13g2_inv_1
X_11469_ _01075_ _05063_ _05045_ VPWR VGND _05064_ sg13g2_nor3_1
X_11470_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _05026_ _05064_ VPWR VGND _00598_ sg13g2_mux2_1
X_11471_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _05013_ _05064_ VPWR VGND _00599_ sg13g2_mux2_1
X_11472_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _05025_ _05064_ VPWR VGND _00600_ sg13g2_mux2_1
X_11473_ _00115_ _05017_ _05064_ VPWR VGND _00601_ sg13g2_mux2_1
X_11474_ _01075_ _05063_ VPWR VGND _05065_ sg13g2_nor2_1
X_11475_ _05034_ _05065_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[6]\ VPWR VGND _05066_ sg13g2_a21oi_1
X_11476_ _05019_ _05065_ _05066_ VPWR VGND _00602_ sg13g2_a21oi_1
X_11477_ _01035_ _01073_ VPWR VGND _05067_ sg13g2_nor2_1
X_11478_ _01068_ _05067_ idle_led_o VPWR VGND _05068_ sg13g2_a21oi_1
X_11479_ _00853_ \atbs_core_0.enable_analog_uart\ _01033_ VPWR VGND _05069_ sg13g2_a21oi_1
X_11480_ _01069_ _04985_ _00845_ _05069_ VPWR VGND 
+ _05070_
+ sg13g2_nor4_1
X_11481_ _05068_ _05070_ VPWR VGND _00603_ sg13g2_nor2_1
X_11482_ _00843_ _00027_ _04982_ VPWR VGND _05071_ sg13g2_nand3_1
X_11483_ overflow_led_o _05071_ _04987_ VPWR VGND _00604_ sg13g2_a21o_1
X_11484_ _05071_ VPWR VGND _05072_ sg13g2_inv_1
X_11485_ _01069_ _04985_ _00843_ _04984_ VPWR VGND 
+ _05073_
+ sg13g2_nand4_1
X_11486_ _00989_ VPWR VGND _05074_ sg13g2_inv_1
X_11487_ _05074_ _04986_ VPWR VGND _05075_ sg13g2_nor2_1
X_11488_ underflow_led_o _05073_ _05075_ VPWR VGND _05076_ sg13g2_a21oi_1
X_11489_ _05072_ _05076_ VPWR VGND _00605_ sg13g2_nor2_1
X_11490_ _01051_ _01053_ VPWR VGND _05077_ sg13g2_nor2_1
X_11491_ \atbs_core_0.atbs_max_delta_steps_uart\ _05063_ _01058_ VPWR VGND _05078_ sg13g2_nor3_1
X_11492_ _01052_ _05077_ _05078_ VPWR VGND _05079_ sg13g2_nand3b_1
X_11493_ _01087_ _00116_ _05079_ VPWR VGND _00606_ sg13g2_mux2_1
X_11494_ _01083_ _05078_ VPWR VGND _05080_ sg13g2_nand2b_1
X_11495_ \atbs_core_0.adaptive_mode_uart\ _05080_ VPWR VGND _05081_ sg13g2_nand2_1
X_11496_ _01087_ _05080_ _05081_ VPWR VGND _00607_ sg13g2_o21ai_1
X_11497_ _05030_ _05078_ VPWR VGND _05082_ sg13g2_nand2_1
X_11498_ _00117_ _05082_ VPWR VGND _05083_ sg13g2_nand2_1
X_11499_ _01048_ _05082_ _05083_ VPWR VGND _00608_ sg13g2_o21ai_1
X_11500_ _01052_ _05077_ _05078_ VPWR VGND _05084_ sg13g2_nand3_1
X_11501_ _00118_ _05084_ VPWR VGND _05085_ sg13g2_nand2_1
X_11502_ _01048_ _05084_ _05085_ VPWR VGND _00609_ sg13g2_o21ai_1
X_11503_ _00944_ _01102_ VPWR VGND _05086_ sg13g2_nor2_1
X_11504_ \atbs_core_0.spike_detector_0.lock_detection\ _05086_ VPWR VGND _05087_ sg13g2_nor2_1
X_11505_ \atbs_core_0.spike_detector_0.is_changing\ _00991_ _05087_ _02109_ VPWR VGND 
+ _00610_
+ sg13g2_a22oi_1
X_11506_ \atbs_core_0.dac_control_0.dac_change_in_progress\ VPWR VGND _05088_ sg13g2_inv_1
X_11507_ _05088_ _04621_ \atbs_core_0.spike_detector_0.n1258_q\ VPWR VGND _05089_ sg13g2_o21ai_1
X_11508_ _00951_ _05089_ VPWR VGND _00611_ sg13g2_nand2_1
X_11509_ \atbs_core_0.dac_control_1.dac_change_in_progress\ VPWR VGND _05090_ sg13g2_inv_1
X_11510_ _05090_ _04829_ \atbs_core_0.spike_detector_0.lower_is_changing\ VPWR VGND _05091_ sg13g2_o21ai_1
X_11511_ _01031_ _05091_ VPWR VGND _00612_ sg13g2_nand2_1
X_11512_ _01097_ \atbs_core_0.spike_encoder_0.delayed_spike_strb\ _01105_ VPWR VGND _05092_ sg13g2_nor3_1
X_11513_ _05092_ VPWR VGND _05093_ sg13g2_buf_1
X_11514_ _05093_ VPWR VGND \atbs_core_0.spike_encoder_0.n1860_o\ sg13g2_inv_1
X_11515_ _05093_ VPWR VGND _05094_ sg13g2_buf_1
X_11516_ _01097_ _01970_ VPWR VGND _05095_ sg13g2_nand2b_1
X_11517_ \atbs_core_0.encoded_spike[0]\ _05094_ VPWR VGND _05096_ sg13g2_nand2_1
X_11518_ _05094_ _05095_ _05096_ VPWR VGND _00613_ sg13g2_o21ai_1
X_11519_ \atbs_core_0.spike_encoder_0.delayed_spike\ \atbs_core_0.adaptive_ctrl_0.spike_i\ VPWR VGND _05097_ sg13g2_nor2_1
X_11520_ _05097_ VPWR VGND _05098_ sg13g2_buf_1
X_11521_ _05098_ VPWR VGND _05099_ sg13g2_buf_1
X_11522_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[9]\ VPWR VGND _05100_ sg13g2_buf_1
X_11523_ _05100_ VPWR VGND _05101_ sg13g2_inv_1
X_11524_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[7]\ VPWR VGND _05102_ sg13g2_buf_1
X_11525_ _01803_ _01810_ _01784_ VPWR VGND _05103_ sg13g2_nor3_1
X_11526_ _01966_ _01972_ _05103_ VPWR VGND _05104_ sg13g2_nand3_1
X_11527_ _01827_ _05102_ _05104_ VPWR VGND _05105_ sg13g2_nor3_1
X_11528_ _04239_ _05105_ VPWR VGND _05106_ sg13g2_and2_1
X_11529_ _05106_ VPWR VGND _05107_ sg13g2_buf_1
X_11530_ _05101_ _05107_ VPWR VGND _05108_ sg13g2_and2_1
X_11531_ _02250_ _05108_ VPWR VGND _05109_ sg13g2_xnor2_1
X_11532_ _02197_ _05098_ VPWR VGND _05110_ sg13g2_nor2_1
X_11533_ _05099_ _05109_ _05110_ VPWR VGND _05111_ sg13g2_a21oi_1
X_11534_ _01103_ \atbs_core_0.spike_encoder_0.n1860_o\ VPWR VGND _05112_ sg13g2_nand2_1
X_11535_ _05112_ VPWR VGND _05113_ sg13g2_buf_1
X_11536_ _05113_ VPWR VGND _05114_ sg13g2_buf_1
X_11537_ \atbs_core_0.encoded_spike[10]\ _05094_ VPWR VGND _05115_ sg13g2_nand2_1
X_11538_ _05111_ _05114_ _05115_ VPWR VGND _00614_ sg13g2_o21ai_1
X_11539_ _05098_ VPWR VGND _05116_ sg13g2_buf_1
X_11540_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[11]\ VPWR VGND _05117_ sg13g2_buf_1
X_11541_ _00061_ VPWR VGND _05118_ sg13g2_inv_1
X_11542_ _01795_ _02382_ _05118_ VPWR VGND _05119_ sg13g2_nor3_1
X_11543_ _05103_ _05119_ VPWR VGND _05120_ sg13g2_nand2_1
X_11544_ _01998_ _01827_ _05102_ _05120_ VPWR VGND 
+ _05121_
+ sg13g2_nor4_1
X_11545_ _01728_ _05101_ _05121_ VPWR VGND _05122_ sg13g2_nand3_1
X_11546_ _05117_ _05122_ VPWR VGND _05123_ sg13g2_xor2_1
X_11547_ _05098_ VPWR VGND _05124_ sg13g2_buf_1
X_11548_ _02731_ _05124_ VPWR VGND _05125_ sg13g2_nor2_1
X_11549_ _05116_ _05123_ _05125_ VPWR VGND _05126_ sg13g2_a21oi_1
X_11550_ \atbs_core_0.encoded_spike[11]\ _05094_ VPWR VGND _05127_ sg13g2_nand2_1
X_11551_ _05114_ _05126_ _05127_ VPWR VGND _00615_ sg13g2_o21ai_1
X_11552_ _02250_ _05100_ _05117_ VPWR VGND _05128_ sg13g2_nor3_1
X_11553_ _05107_ _05128_ VPWR VGND _05129_ sg13g2_nand2_1
X_11554_ _02572_ _05129_ VPWR VGND _05130_ sg13g2_xnor2_1
X_11555_ _01856_ _05124_ VPWR VGND _05131_ sg13g2_nor2_1
X_11556_ _05116_ _05130_ _05131_ VPWR VGND _05132_ sg13g2_a21oi_1
X_11557_ \atbs_core_0.encoded_spike[12]\ _05094_ VPWR VGND _05133_ sg13g2_nand2_1
X_11558_ _05114_ _05132_ _05133_ VPWR VGND _00616_ sg13g2_o21ai_1
X_11559_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[13]\ VPWR VGND _05134_ sg13g2_inv_1
X_11560_ _02572_ _05128_ VPWR VGND _05135_ sg13g2_and2_1
X_11561_ _05121_ _05135_ VPWR VGND _05136_ sg13g2_nand2_1
X_11562_ _05134_ _05136_ VPWR VGND _05137_ sg13g2_xnor2_1
X_11563_ _02575_ _05124_ VPWR VGND _05138_ sg13g2_nor2_1
X_11564_ _05116_ _05137_ _05138_ VPWR VGND _05139_ sg13g2_a21oi_1
X_11565_ \atbs_core_0.encoded_spike[13]\ _05094_ VPWR VGND _05140_ sg13g2_nand2_1
X_11566_ _05114_ _05139_ _05140_ VPWR VGND _00617_ sg13g2_o21ai_1
X_11567_ _05134_ _05135_ VPWR VGND _05141_ sg13g2_and2_1
X_11568_ _05107_ _05141_ VPWR VGND _05142_ sg13g2_nand2_1
X_11569_ _01703_ _05142_ VPWR VGND _05143_ sg13g2_xnor2_1
X_11570_ _02428_ _05124_ VPWR VGND _05144_ sg13g2_nor2_1
X_11571_ _05116_ _05143_ _05144_ VPWR VGND _05145_ sg13g2_a21oi_1
X_11572_ \atbs_core_0.encoded_spike[14]\ _05094_ VPWR VGND _05146_ sg13g2_nand2_1
X_11573_ _05114_ _05145_ _05146_ VPWR VGND _00618_ sg13g2_o21ai_1
X_11574_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[15]\ VPWR VGND _05147_ sg13g2_buf_1
X_11575_ _01703_ _05141_ VPWR VGND _05148_ sg13g2_and2_1
X_11576_ _05121_ _05148_ VPWR VGND _05149_ sg13g2_nand2_1
X_11577_ _05147_ _05149_ VPWR VGND _05150_ sg13g2_xor2_1
X_11578_ _02276_ _05124_ VPWR VGND _05151_ sg13g2_nor2_1
X_11579_ _05116_ _05150_ _05151_ VPWR VGND _05152_ sg13g2_a21oi_1
X_11580_ \atbs_core_0.encoded_spike[15]\ _05094_ VPWR VGND _05153_ sg13g2_nand2_1
X_11581_ _05114_ _05152_ _05153_ VPWR VGND _00619_ sg13g2_o21ai_1
X_11582_ _05147_ _05148_ VPWR VGND _05154_ sg13g2_nor2b_1
X_11583_ _05107_ _05154_ VPWR VGND _05155_ sg13g2_nand2_1
X_11584_ _03396_ _05155_ VPWR VGND _05156_ sg13g2_xnor2_1
X_11585_ _02278_ _05124_ VPWR VGND _05157_ sg13g2_nor2_1
X_11586_ _05116_ _05156_ _05157_ VPWR VGND _05158_ sg13g2_a21oi_1
X_11587_ \atbs_core_0.encoded_spike[16]\ _05094_ VPWR VGND _05159_ sg13g2_nand2_1
X_11588_ _05114_ _05158_ _05159_ VPWR VGND _00620_ sg13g2_o21ai_1
X_11589_ _03396_ _05121_ _05154_ VPWR VGND _05160_ sg13g2_nand3_1
X_11590_ _01895_ _05160_ VPWR VGND _05161_ sg13g2_xnor2_1
X_11591_ _01897_ _05124_ VPWR VGND _05162_ sg13g2_nor2_1
X_11592_ _05116_ _05161_ _05162_ VPWR VGND _05163_ sg13g2_a21oi_1
X_11593_ _05093_ VPWR VGND _05164_ sg13g2_buf_1
X_11594_ \atbs_core_0.encoded_spike[17]\ _05164_ VPWR VGND _05165_ sg13g2_nand2_1
X_11595_ _05114_ _05163_ _05165_ VPWR VGND _00621_ sg13g2_o21ai_1
X_11596_ _01895_ _03396_ _05107_ _05154_ VPWR VGND 
+ _05166_
+ sg13g2_nand4_1
X_11597_ _01103_ _05116_ _05166_ VPWR VGND _05167_ sg13g2_nand3_1
X_11598_ \atbs_core_0.encoded_spike[18]\ _05164_ VPWR VGND _05168_ sg13g2_nand2_1
X_11599_ _05094_ _05167_ _05168_ VPWR VGND _00622_ sg13g2_o21ai_1
X_11600_ _01795_ _01970_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[1]\ sg13g2_xor2_1
X_11601_ _00062_ _05124_ VPWR VGND _05169_ sg13g2_nor2_1
X_11602_ _05116_ \atbs_core_0.time_measurement_0.n1813_o[1]\ _05169_ VPWR VGND _05170_ sg13g2_a21oi_1
X_11603_ \atbs_core_0.encoded_spike[1]\ _05164_ VPWR VGND _05171_ sg13g2_nand2_1
X_11604_ _05114_ _05170_ _05171_ VPWR VGND _00623_ sg13g2_o21ai_1
X_11605_ _02382_ _01972_ VPWR VGND _05172_ sg13g2_xnor2_1
X_11606_ _00063_ _05124_ VPWR VGND _05173_ sg13g2_nor2_1
X_11607_ _05116_ _05172_ _05173_ VPWR VGND _05174_ sg13g2_a21oi_1
X_11608_ \atbs_core_0.encoded_spike[2]\ _05164_ VPWR VGND _05175_ sg13g2_nand2_1
X_11609_ _05114_ _05174_ _05175_ VPWR VGND _00624_ sg13g2_o21ai_1
X_11610_ _01803_ _05119_ VPWR VGND _05176_ sg13g2_xnor2_1
X_11611_ _00064_ _05098_ VPWR VGND _05177_ sg13g2_nor2_1
X_11612_ _05099_ _05176_ _05177_ VPWR VGND _05178_ sg13g2_a21oi_1
X_11613_ \atbs_core_0.encoded_spike[3]\ _05164_ VPWR VGND _05179_ sg13g2_nand2_1
X_11614_ _05113_ _05178_ _05179_ VPWR VGND _00625_ sg13g2_o21ai_1
X_11615_ _01795_ _01970_ _01803_ _02382_ VPWR VGND 
+ _05180_
+ sg13g2_nor4_1
X_11616_ _01784_ _05180_ VPWR VGND _05181_ sg13g2_xnor2_1
X_11617_ _00065_ _05098_ VPWR VGND _05182_ sg13g2_nor2_1
X_11618_ _05099_ _05181_ _05182_ VPWR VGND _05183_ sg13g2_a21oi_1
X_11619_ \atbs_core_0.encoded_spike[4]\ _05164_ VPWR VGND _05184_ sg13g2_nand2_1
X_11620_ _05113_ _05183_ _05184_ VPWR VGND _00626_ sg13g2_o21ai_1
X_11621_ _02222_ _01964_ _05119_ VPWR VGND _05185_ sg13g2_nand3_1
X_11622_ _01980_ _05185_ VPWR VGND _05186_ sg13g2_xnor2_1
X_11623_ _00066_ _05098_ VPWR VGND _05187_ sg13g2_nor2_1
X_11624_ _05099_ _05186_ _05187_ VPWR VGND _05188_ sg13g2_a21oi_1
X_11625_ \atbs_core_0.encoded_spike[5]\ _05164_ VPWR VGND _05189_ sg13g2_nand2_1
X_11626_ _05113_ _05188_ _05189_ VPWR VGND _00627_ sg13g2_o21ai_1
X_11627_ _01827_ _05104_ VPWR VGND _05190_ sg13g2_xnor2_1
X_11628_ _05099_ _05190_ VPWR VGND _05191_ sg13g2_nand2_1
X_11629_ _01962_ _05099_ _05191_ VPWR VGND _05192_ sg13g2_o21ai_1
X_11630_ \atbs_core_0.encoded_spike[6]\ _05164_ VPWR VGND _05193_ sg13g2_nand2_1
X_11631_ _05113_ _05192_ _05193_ VPWR VGND _00628_ sg13g2_o21ai_1
X_11632_ _05102_ VPWR VGND _05194_ sg13g2_inv_1
X_11633_ _01827_ _05120_ VPWR VGND _05195_ sg13g2_nor2_1
X_11634_ _05194_ _05195_ VPWR VGND _05196_ sg13g2_xnor2_1
X_11635_ _05099_ _05196_ VPWR VGND _05197_ sg13g2_nand2_1
X_11636_ _02548_ _05099_ _05197_ VPWR VGND _05198_ sg13g2_o21ai_1
X_11637_ \atbs_core_0.encoded_spike[7]\ _05164_ VPWR VGND _05199_ sg13g2_nand2_1
X_11638_ _05113_ _05198_ _05199_ VPWR VGND _00629_ sg13g2_o21ai_1
X_11639_ _04239_ _05105_ VPWR VGND _05200_ sg13g2_nor2_1
X_11640_ _05107_ _05200_ _05098_ VPWR VGND _05201_ sg13g2_o21ai_1
X_11641_ _01989_ _05099_ _05201_ VPWR VGND _05202_ sg13g2_o21ai_1
X_11642_ \atbs_core_0.encoded_spike[8]\ _05164_ VPWR VGND _05203_ sg13g2_nand2_1
X_11643_ _05113_ _05202_ _05203_ VPWR VGND _00630_ sg13g2_o21ai_1
X_11644_ _05101_ _05121_ VPWR VGND _05204_ sg13g2_xnor2_1
X_11645_ _05124_ _05204_ VPWR VGND _05205_ sg13g2_nand2_1
X_11646_ _02687_ _05099_ _05205_ VPWR VGND _05206_ sg13g2_o21ai_1
X_11647_ \atbs_core_0.encoded_spike[9]\ _05093_ VPWR VGND _05207_ sg13g2_nand2_1
X_11648_ _05113_ _05206_ _05207_ VPWR VGND _00631_ sg13g2_o21ai_1
X_11649_ \atbs_core_0.spike_memory_0.n1974_q\ VPWR VGND _05208_ sg13g2_buf_1
X_11650_ _05208_ VPWR VGND _05209_ sg13g2_buf_1
X_11651_ _05209_ VPWR VGND _05210_ sg13g2_buf_1
X_11652_ \atbs_core_0.spike_memory_0.n1953_o[0]\ \atbs_core_0.spike_memory_0.a_data[0]\ _05210_ VPWR VGND _00632_ sg13g2_mux2_1
X_11653_ \atbs_core_0.spike_memory_0.n1953_o[10]\ \atbs_core_0.spike_memory_0.a_data[10]\ _05210_ VPWR VGND _00633_ sg13g2_mux2_1
X_11654_ \atbs_core_0.spike_memory_0.n1953_o[11]\ \atbs_core_0.spike_memory_0.a_data[11]\ _05210_ VPWR VGND _00634_ sg13g2_mux2_1
X_11655_ \atbs_core_0.spike_memory_0.n1953_o[12]\ \atbs_core_0.spike_memory_0.a_data[12]\ _05210_ VPWR VGND _00635_ sg13g2_mux2_1
X_11656_ \atbs_core_0.spike_memory_0.n1953_o[13]\ \atbs_core_0.spike_memory_0.a_data[13]\ _05210_ VPWR VGND _00636_ sg13g2_mux2_1
X_11657_ \atbs_core_0.spike_memory_0.n1953_o[14]\ \atbs_core_0.spike_memory_0.a_data[14]\ _05210_ VPWR VGND _00637_ sg13g2_mux2_1
X_11658_ \atbs_core_0.spike_memory_0.n1953_o[15]\ \atbs_core_0.spike_memory_0.a_data[15]\ _05210_ VPWR VGND _00638_ sg13g2_mux2_1
X_11659_ \atbs_core_0.spike_memory_0.n1953_o[16]\ \atbs_core_0.spike_memory_0.a_data[16]\ _05210_ VPWR VGND _00639_ sg13g2_mux2_1
X_11660_ \atbs_core_0.spike_memory_0.n1953_o[17]\ \atbs_core_0.spike_memory_0.a_data[17]\ _05210_ VPWR VGND _00640_ sg13g2_mux2_1
X_11661_ \atbs_core_0.spike_memory_0.n1953_o[18]\ \atbs_core_0.spike_memory_0.a_data[18]\ _05210_ VPWR VGND _00641_ sg13g2_mux2_1
X_11662_ _05209_ VPWR VGND _05211_ sg13g2_buf_1
X_11663_ \atbs_core_0.spike_memory_0.n1954_o[0]\ \atbs_core_0.spike_memory_0.n1953_o[0]\ _05211_ VPWR VGND _00642_ sg13g2_mux2_1
X_11664_ \atbs_core_0.spike_memory_0.n1953_o[1]\ \atbs_core_0.spike_memory_0.a_data[1]\ _05211_ VPWR VGND _00643_ sg13g2_mux2_1
X_11665_ \atbs_core_0.spike_memory_0.n1954_o[1]\ \atbs_core_0.spike_memory_0.n1953_o[1]\ _05211_ VPWR VGND _00644_ sg13g2_mux2_1
X_11666_ \atbs_core_0.spike_memory_0.n1954_o[2]\ \atbs_core_0.spike_memory_0.n1953_o[2]\ _05211_ VPWR VGND _00645_ sg13g2_mux2_1
X_11667_ \atbs_core_0.spike_memory_0.n1954_o[3]\ \atbs_core_0.spike_memory_0.n1953_o[3]\ _05211_ VPWR VGND _00646_ sg13g2_mux2_1
X_11668_ \atbs_core_0.spike_memory_0.n1954_o[4]\ \atbs_core_0.spike_memory_0.n1953_o[4]\ _05211_ VPWR VGND _00647_ sg13g2_mux2_1
X_11669_ \atbs_core_0.spike_memory_0.n1954_o[5]\ \atbs_core_0.spike_memory_0.n1953_o[5]\ _05211_ VPWR VGND _00648_ sg13g2_mux2_1
X_11670_ \atbs_core_0.spike_memory_0.n1954_o[6]\ \atbs_core_0.spike_memory_0.n1953_o[6]\ _05211_ VPWR VGND _00649_ sg13g2_mux2_1
X_11671_ \atbs_core_0.spike_memory_0.n1954_o[7]\ \atbs_core_0.spike_memory_0.n1953_o[7]\ _05211_ VPWR VGND _00650_ sg13g2_mux2_1
X_11672_ \atbs_core_0.spike_memory_0.n1954_o[8]\ \atbs_core_0.spike_memory_0.n1953_o[8]\ _05211_ VPWR VGND _00651_ sg13g2_mux2_1
X_11673_ _05209_ VPWR VGND _05212_ sg13g2_buf_1
X_11674_ \atbs_core_0.spike_memory_0.n1954_o[9]\ \atbs_core_0.spike_memory_0.n1953_o[9]\ _05212_ VPWR VGND _00652_ sg13g2_mux2_1
X_11675_ \atbs_core_0.spike_memory_0.n1954_o[10]\ \atbs_core_0.spike_memory_0.n1953_o[10]\ _05212_ VPWR VGND _00653_ sg13g2_mux2_1
X_11676_ \atbs_core_0.spike_memory_0.n1953_o[2]\ \atbs_core_0.spike_memory_0.a_data[2]\ _05212_ VPWR VGND _00654_ sg13g2_mux2_1
X_11677_ \atbs_core_0.spike_memory_0.n1954_o[11]\ \atbs_core_0.spike_memory_0.n1953_o[11]\ _05212_ VPWR VGND _00655_ sg13g2_mux2_1
X_11678_ \atbs_core_0.spike_memory_0.n1954_o[12]\ \atbs_core_0.spike_memory_0.n1953_o[12]\ _05212_ VPWR VGND _00656_ sg13g2_mux2_1
X_11679_ \atbs_core_0.spike_memory_0.n1954_o[13]\ \atbs_core_0.spike_memory_0.n1953_o[13]\ _05212_ VPWR VGND _00657_ sg13g2_mux2_1
X_11680_ \atbs_core_0.spike_memory_0.n1954_o[14]\ \atbs_core_0.spike_memory_0.n1953_o[14]\ _05212_ VPWR VGND _00658_ sg13g2_mux2_1
X_11681_ \atbs_core_0.spike_memory_0.n1954_o[15]\ \atbs_core_0.spike_memory_0.n1953_o[15]\ _05212_ VPWR VGND _00659_ sg13g2_mux2_1
X_11682_ \atbs_core_0.spike_memory_0.n1954_o[16]\ \atbs_core_0.spike_memory_0.n1953_o[16]\ _05212_ VPWR VGND _00660_ sg13g2_mux2_1
X_11683_ \atbs_core_0.spike_memory_0.n1954_o[17]\ \atbs_core_0.spike_memory_0.n1953_o[17]\ _05212_ VPWR VGND _00661_ sg13g2_mux2_1
X_11684_ _05209_ VPWR VGND _05213_ sg13g2_buf_1
X_11685_ \atbs_core_0.spike_memory_0.n1954_o[18]\ \atbs_core_0.spike_memory_0.n1953_o[18]\ _05213_ VPWR VGND _00662_ sg13g2_mux2_1
X_11686_ \atbs_core_0.spike_memory_0.n1955_o[0]\ \atbs_core_0.spike_memory_0.n1954_o[0]\ _05213_ VPWR VGND _00663_ sg13g2_mux2_1
X_11687_ \atbs_core_0.spike_memory_0.n1955_o[1]\ \atbs_core_0.spike_memory_0.n1954_o[1]\ _05213_ VPWR VGND _00664_ sg13g2_mux2_1
X_11688_ \atbs_core_0.spike_memory_0.n1953_o[3]\ \atbs_core_0.spike_memory_0.a_data[3]\ _05213_ VPWR VGND _00665_ sg13g2_mux2_1
X_11689_ \atbs_core_0.spike_memory_0.n1955_o[2]\ \atbs_core_0.spike_memory_0.n1954_o[2]\ _05213_ VPWR VGND _00666_ sg13g2_mux2_1
X_11690_ \atbs_core_0.spike_memory_0.n1955_o[3]\ \atbs_core_0.spike_memory_0.n1954_o[3]\ _05213_ VPWR VGND _00667_ sg13g2_mux2_1
X_11691_ \atbs_core_0.spike_memory_0.n1955_o[4]\ \atbs_core_0.spike_memory_0.n1954_o[4]\ _05213_ VPWR VGND _00668_ sg13g2_mux2_1
X_11692_ \atbs_core_0.spike_memory_0.n1955_o[5]\ \atbs_core_0.spike_memory_0.n1954_o[5]\ _05213_ VPWR VGND _00669_ sg13g2_mux2_1
X_11693_ \atbs_core_0.spike_memory_0.n1955_o[6]\ \atbs_core_0.spike_memory_0.n1954_o[6]\ _05213_ VPWR VGND _00670_ sg13g2_mux2_1
X_11694_ \atbs_core_0.spike_memory_0.n1955_o[7]\ \atbs_core_0.spike_memory_0.n1954_o[7]\ _05213_ VPWR VGND _00671_ sg13g2_mux2_1
X_11695_ _05208_ VPWR VGND _05214_ sg13g2_buf_1
X_11696_ \atbs_core_0.spike_memory_0.n1955_o[8]\ \atbs_core_0.spike_memory_0.n1954_o[8]\ _05214_ VPWR VGND _00672_ sg13g2_mux2_1
X_11697_ \atbs_core_0.spike_memory_0.n1955_o[9]\ \atbs_core_0.spike_memory_0.n1954_o[9]\ _05214_ VPWR VGND _00673_ sg13g2_mux2_1
X_11698_ \atbs_core_0.spike_memory_0.n1955_o[10]\ \atbs_core_0.spike_memory_0.n1954_o[10]\ _05214_ VPWR VGND _00674_ sg13g2_mux2_1
X_11699_ \atbs_core_0.spike_memory_0.n1955_o[11]\ \atbs_core_0.spike_memory_0.n1954_o[11]\ _05214_ VPWR VGND _00675_ sg13g2_mux2_1
X_11700_ \atbs_core_0.spike_memory_0.n1953_o[4]\ \atbs_core_0.spike_memory_0.a_data[4]\ _05214_ VPWR VGND _00676_ sg13g2_mux2_1
X_11701_ \atbs_core_0.spike_memory_0.n1955_o[12]\ \atbs_core_0.spike_memory_0.n1954_o[12]\ _05214_ VPWR VGND _00677_ sg13g2_mux2_1
X_11702_ \atbs_core_0.spike_memory_0.n1955_o[13]\ \atbs_core_0.spike_memory_0.n1954_o[13]\ _05214_ VPWR VGND _00678_ sg13g2_mux2_1
X_11703_ \atbs_core_0.spike_memory_0.n1955_o[14]\ \atbs_core_0.spike_memory_0.n1954_o[14]\ _05214_ VPWR VGND _00679_ sg13g2_mux2_1
X_11704_ \atbs_core_0.spike_memory_0.n1955_o[15]\ \atbs_core_0.spike_memory_0.n1954_o[15]\ _05214_ VPWR VGND _00680_ sg13g2_mux2_1
X_11705_ \atbs_core_0.spike_memory_0.n1955_o[16]\ \atbs_core_0.spike_memory_0.n1954_o[16]\ _05214_ VPWR VGND _00681_ sg13g2_mux2_1
X_11706_ _05208_ VPWR VGND _05215_ sg13g2_buf_1
X_11707_ \atbs_core_0.spike_memory_0.n1955_o[17]\ \atbs_core_0.spike_memory_0.n1954_o[17]\ _05215_ VPWR VGND _00682_ sg13g2_mux2_1
X_11708_ \atbs_core_0.spike_memory_0.n1955_o[18]\ \atbs_core_0.spike_memory_0.n1954_o[18]\ _05215_ VPWR VGND _00683_ sg13g2_mux2_1
X_11709_ \atbs_core_0.spike_memory_0.n1971_q[57]\ \atbs_core_0.spike_memory_0.n1955_o[0]\ _05215_ VPWR VGND _00684_ sg13g2_mux2_1
X_11710_ \atbs_core_0.spike_memory_0.n1971_q[58]\ \atbs_core_0.spike_memory_0.n1955_o[1]\ _05215_ VPWR VGND _00685_ sg13g2_mux2_1
X_11711_ \atbs_core_0.spike_memory_0.n1971_q[59]\ \atbs_core_0.spike_memory_0.n1955_o[2]\ _05215_ VPWR VGND _00686_ sg13g2_mux2_1
X_11712_ \atbs_core_0.spike_memory_0.n1953_o[5]\ \atbs_core_0.spike_memory_0.a_data[5]\ _05215_ VPWR VGND _00687_ sg13g2_mux2_1
X_11713_ \atbs_core_0.spike_memory_0.n1971_q[60]\ \atbs_core_0.spike_memory_0.n1955_o[3]\ _05215_ VPWR VGND _00688_ sg13g2_mux2_1
X_11714_ \atbs_core_0.spike_memory_0.n1971_q[61]\ \atbs_core_0.spike_memory_0.n1955_o[4]\ _05215_ VPWR VGND _00689_ sg13g2_mux2_1
X_11715_ \atbs_core_0.spike_memory_0.n1971_q[62]\ \atbs_core_0.spike_memory_0.n1955_o[5]\ _05215_ VPWR VGND _00690_ sg13g2_mux2_1
X_11716_ \atbs_core_0.spike_memory_0.n1971_q[63]\ \atbs_core_0.spike_memory_0.n1955_o[6]\ _05215_ VPWR VGND _00691_ sg13g2_mux2_1
X_11717_ _05208_ VPWR VGND _05216_ sg13g2_buf_1
X_11718_ \atbs_core_0.spike_memory_0.n1971_q[64]\ \atbs_core_0.spike_memory_0.n1955_o[7]\ _05216_ VPWR VGND _00692_ sg13g2_mux2_1
X_11719_ \atbs_core_0.spike_memory_0.n1971_q[65]\ \atbs_core_0.spike_memory_0.n1955_o[8]\ _05216_ VPWR VGND _00693_ sg13g2_mux2_1
X_11720_ \atbs_core_0.spike_memory_0.n1971_q[66]\ \atbs_core_0.spike_memory_0.n1955_o[9]\ _05216_ VPWR VGND _00694_ sg13g2_mux2_1
X_11721_ \atbs_core_0.spike_memory_0.n1971_q[67]\ \atbs_core_0.spike_memory_0.n1955_o[10]\ _05216_ VPWR VGND _00695_ sg13g2_mux2_1
X_11722_ \atbs_core_0.spike_memory_0.n1971_q[68]\ \atbs_core_0.spike_memory_0.n1955_o[11]\ _05216_ VPWR VGND _00696_ sg13g2_mux2_1
X_11723_ \atbs_core_0.spike_memory_0.n1971_q[69]\ \atbs_core_0.spike_memory_0.n1955_o[12]\ _05216_ VPWR VGND _00697_ sg13g2_mux2_1
X_11724_ \atbs_core_0.spike_memory_0.n1953_o[6]\ \atbs_core_0.spike_memory_0.a_data[6]\ _05216_ VPWR VGND _00698_ sg13g2_mux2_1
X_11725_ \atbs_core_0.spike_memory_0.n1971_q[70]\ \atbs_core_0.spike_memory_0.n1955_o[13]\ _05216_ VPWR VGND _00699_ sg13g2_mux2_1
X_11726_ \atbs_core_0.spike_memory_0.n1971_q[71]\ \atbs_core_0.spike_memory_0.n1955_o[14]\ _05216_ VPWR VGND _00700_ sg13g2_mux2_1
X_11727_ \atbs_core_0.spike_memory_0.n1971_q[72]\ \atbs_core_0.spike_memory_0.n1955_o[15]\ _05216_ VPWR VGND _00701_ sg13g2_mux2_1
X_11728_ \atbs_core_0.spike_memory_0.n1971_q[73]\ \atbs_core_0.spike_memory_0.n1955_o[16]\ _05209_ VPWR VGND _00702_ sg13g2_mux2_1
X_11729_ \atbs_core_0.spike_memory_0.n1971_q[74]\ \atbs_core_0.spike_memory_0.n1955_o[17]\ _05209_ VPWR VGND _00703_ sg13g2_mux2_1
X_11730_ \atbs_core_0.spike_memory_0.n1971_q[75]\ \atbs_core_0.spike_memory_0.n1955_o[18]\ _05209_ VPWR VGND _00704_ sg13g2_mux2_1
X_11731_ \atbs_core_0.spike_memory_0.n1953_o[7]\ \atbs_core_0.spike_memory_0.a_data[7]\ _05209_ VPWR VGND _00705_ sg13g2_mux2_1
X_11732_ \atbs_core_0.spike_memory_0.n1953_o[8]\ \atbs_core_0.spike_memory_0.a_data[8]\ _05209_ VPWR VGND _00706_ sg13g2_mux2_1
X_11733_ \atbs_core_0.spike_memory_0.n1953_o[9]\ \atbs_core_0.spike_memory_0.a_data[9]\ _05209_ VPWR VGND _00707_ sg13g2_mux2_1
X_11734_ \atbs_core_0.encoded_spike_strb\ \atbs_core_0.n1056_q\ _04984_ VPWR VGND _05217_ sg13g2_and3_1
X_11735_ _05217_ VPWR VGND _05218_ sg13g2_buf_1
X_11736_ _05218_ VPWR VGND \atbs_core_0.spike_memory_0.n1899_o\ sg13g2_buf_1
X_11737_ _00986_ VPWR VGND _05219_ sg13g2_buf_1
X_11738_ _05219_ VPWR VGND _05220_ sg13g2_buf_1
X_11739_ _05220_ \atbs_core_0.spike_memory_0.n1901_o[0]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00708_ sg13g2_mux2_1
X_11740_ _05220_ _05218_ VPWR VGND _05221_ sg13g2_nand2_1
X_11741_ \atbs_core_0.spike_memory_0.head[1]\ _05221_ VPWR VGND _00709_ sg13g2_xnor2_1
X_11742_ _00985_ VPWR VGND _05222_ sg13g2_buf_1
X_11743_ _05222_ \atbs_core_0.spike_memory_0.n1916_o[0]\ \atbs_core_0.spike_memory_0.n1914_o\ VPWR VGND _00710_ sg13g2_mux2_1
X_11744_ _05222_ \atbs_core_0.spike_memory_0.n1914_o\ VPWR VGND _05223_ sg13g2_nand2_1
X_11745_ \atbs_core_0.spike_memory_0.n1973_q[1]\ _05223_ VPWR VGND _00711_ sg13g2_xnor2_1
X_11746_ \atbs_core_0.spike_memory_0.a_data[0]\ \atbs_core_0.encoded_spike[0]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00712_ sg13g2_mux2_1
X_11747_ \atbs_core_0.spike_memory_0.a_data[10]\ \atbs_core_0.encoded_spike[10]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00713_ sg13g2_mux2_1
X_11748_ \atbs_core_0.spike_memory_0.a_data[11]\ \atbs_core_0.encoded_spike[11]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00714_ sg13g2_mux2_1
X_11749_ \atbs_core_0.spike_memory_0.a_data[12]\ \atbs_core_0.encoded_spike[12]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00715_ sg13g2_mux2_1
X_11750_ \atbs_core_0.spike_memory_0.a_data[13]\ \atbs_core_0.encoded_spike[13]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00716_ sg13g2_mux2_1
X_11751_ \atbs_core_0.spike_memory_0.a_data[14]\ \atbs_core_0.encoded_spike[14]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00717_ sg13g2_mux2_1
X_11752_ \atbs_core_0.spike_memory_0.a_data[15]\ \atbs_core_0.encoded_spike[15]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00718_ sg13g2_mux2_1
X_11753_ \atbs_core_0.spike_memory_0.a_data[16]\ \atbs_core_0.encoded_spike[16]\ \atbs_core_0.spike_memory_0.n1899_o\ VPWR VGND _00719_ sg13g2_mux2_1
X_11754_ _05218_ VPWR VGND _05224_ sg13g2_buf_1
X_11755_ \atbs_core_0.spike_memory_0.a_data[17]\ \atbs_core_0.encoded_spike[17]\ _05224_ VPWR VGND _00720_ sg13g2_mux2_1
X_11756_ \atbs_core_0.spike_memory_0.a_data[18]\ \atbs_core_0.encoded_spike[18]\ _05224_ VPWR VGND _00721_ sg13g2_mux2_1
X_11757_ \atbs_core_0.spike_memory_0.a_data[1]\ \atbs_core_0.encoded_spike[1]\ _05224_ VPWR VGND _00722_ sg13g2_mux2_1
X_11758_ \atbs_core_0.spike_memory_0.a_data[2]\ \atbs_core_0.encoded_spike[2]\ _05224_ VPWR VGND _00723_ sg13g2_mux2_1
X_11759_ \atbs_core_0.spike_memory_0.a_data[3]\ \atbs_core_0.encoded_spike[3]\ _05224_ VPWR VGND _00724_ sg13g2_mux2_1
X_11760_ \atbs_core_0.spike_memory_0.a_data[4]\ \atbs_core_0.encoded_spike[4]\ _05224_ VPWR VGND _00725_ sg13g2_mux2_1
X_11761_ \atbs_core_0.spike_memory_0.a_data[5]\ \atbs_core_0.encoded_spike[5]\ _05224_ VPWR VGND _00726_ sg13g2_mux2_1
X_11762_ \atbs_core_0.spike_memory_0.a_data[6]\ \atbs_core_0.encoded_spike[6]\ _05224_ VPWR VGND _00727_ sg13g2_mux2_1
X_11763_ \atbs_core_0.spike_memory_0.a_data[7]\ \atbs_core_0.encoded_spike[7]\ _05224_ VPWR VGND _00728_ sg13g2_mux2_1
X_11764_ \atbs_core_0.spike_memory_0.a_data[8]\ \atbs_core_0.encoded_spike[8]\ _05224_ VPWR VGND _00729_ sg13g2_mux2_1
X_11765_ \atbs_core_0.spike_memory_0.a_data[9]\ \atbs_core_0.encoded_spike[9]\ _05218_ VPWR VGND _00730_ sg13g2_mux2_1
X_11766_ \atbs_core_0.memory2uart_0.tx_strb_i\ \atbs_core_0.spike_memory_0.n1914_o\ VPWR VGND _05225_ sg13g2_nor2_1
X_11767_ \atbs_core_0.spike_memory_0.n1928_o[0]\ \atbs_core_0.spike_memory_0.n1926_o\ _05225_ VPWR VGND _00731_ sg13g2_mux2_1
X_11768_ \atbs_core_0.spike_memory_0.n1926_o\ VPWR VGND _05226_ sg13g2_inv_1
X_11769_ \atbs_core_0.spike_memory_0.n1925_o\ \atbs_core_0.spike_memory_0.n1914_o\ _04926_ VPWR VGND _05227_ sg13g2_o21ai_1
X_11770_ _04926_ _05226_ _05227_ VPWR VGND _00732_ sg13g2_o21ai_1
X_11771_ \atbs_core_0.spike_memory_0.n1925_o\ VPWR VGND _05228_ sg13g2_inv_1
X_11772_ \atbs_core_0.spike_memory_0.n1912_o\ \atbs_core_0.spike_memory_0.n1914_o\ _04926_ VPWR VGND _05229_ sg13g2_o21ai_1
X_11773_ _04926_ _05228_ _05229_ VPWR VGND _00733_ sg13g2_o21ai_1
X_11774_ _00787_ _00784_ VPWR VGND _05230_ sg13g2_xnor2_1
X_11775_ _00789_ _05230_ VPWR VGND _00734_ sg13g2_and2_1
X_11776_ _00785_ _00954_ VPWR VGND _05231_ sg13g2_xnor2_1
X_11777_ _00789_ _05231_ VPWR VGND _00735_ sg13g2_and2_1
X_11778_ _00785_ _00787_ _00953_ VPWR VGND _05232_ sg13g2_nand3_1
X_11779_ _00786_ _05232_ VPWR VGND _05233_ sg13g2_xnor2_1
X_11780_ _00789_ _05233_ VPWR VGND _00736_ sg13g2_and2_1
X_11781_ _00785_ _00786_ VPWR VGND _05234_ sg13g2_nor2_1
X_11782_ _00007_ _05234_ VPWR VGND _05235_ sg13g2_nand2_1
X_11783_ _00961_ _00964_ _00968_ VPWR VGND _05236_ sg13g2_nand3b_1
X_11784_ _00956_ _00789_ VPWR VGND _05237_ sg13g2_nand2b_1
X_11785_ _00748_ _00971_ _05236_ _05237_ VPWR VGND 
+ _05238_
+ sg13g2_nor4_1
X_11786_ _05238_ VPWR VGND _05239_ sg13g2_buf_1
X_11787_ _00789_ _00956_ VPWR VGND _05240_ sg13g2_nor2_1
X_11788_ _00789_ _00956_ VPWR VGND _05241_ sg13g2_nand2b_1
X_11789_ _05237_ _00969_ VPWR VGND _05242_ sg13g2_nand2b_1
X_11790_ _05241_ _05242_ _00971_ VPWR VGND _05243_ sg13g2_a21oi_1
X_11791_ _00971_ _05240_ _05243_ VPWR VGND _05244_ sg13g2_a21oi_1
X_11792_ _00971_ _05240_ _00748_ VPWR VGND _05245_ sg13g2_nand3b_1
X_11793_ _00748_ _05244_ _05245_ VPWR VGND _05246_ sg13g2_o21ai_1
X_11794_ _05246_ VPWR VGND _05247_ sg13g2_buf_1
X_11795_ _05235_ _05239_ _05247_ VPWR VGND _05248_ sg13g2_a21oi_1
X_11796_ _00748_ _00971_ _00972_ _05237_ VPWR VGND 
+ _05249_
+ sg13g2_nor4_1
X_11797_ _05249_ VPWR VGND _05250_ sg13g2_buf_1
X_11798_ _05250_ _05248_ VPWR VGND _05251_ sg13g2_nand2_1
X_11799_ _01087_ _05248_ _05251_ VPWR VGND _00737_ sg13g2_o21ai_1
X_11800_ _00787_ _05234_ VPWR VGND _05252_ sg13g2_nand2_1
X_11801_ _05239_ _05252_ _05247_ VPWR VGND _05253_ sg13g2_a21oi_1
X_11802_ _01051_ _05250_ _05253_ VPWR VGND _00738_ sg13g2_mux2_1
X_11803_ _00786_ _00007_ _00785_ VPWR VGND _05254_ sg13g2_nand3b_1
X_11804_ _05239_ _05254_ _05247_ VPWR VGND _05255_ sg13g2_a21oi_1
X_11805_ _01053_ _05250_ _05255_ VPWR VGND _00739_ sg13g2_mux2_1
X_11806_ _00786_ _00787_ _00785_ VPWR VGND _05256_ sg13g2_nand3b_1
X_11807_ _05239_ _05256_ _05247_ VPWR VGND _05257_ sg13g2_a21oi_1
X_11808_ _01052_ _05250_ _05257_ VPWR VGND _00740_ sg13g2_mux2_1
X_11809_ _00785_ _00786_ _00007_ VPWR VGND _05258_ sg13g2_nand3b_1
X_11810_ _05239_ _05258_ _05247_ VPWR VGND _05259_ sg13g2_a21oi_1
X_11811_ _05250_ _05259_ VPWR VGND _05260_ sg13g2_nand2_1
X_11812_ _01044_ _05259_ _05260_ VPWR VGND _00741_ sg13g2_o21ai_1
X_11813_ _00785_ _00786_ _00787_ VPWR VGND _05261_ sg13g2_nand3b_1
X_11814_ _05239_ _05261_ _05247_ VPWR VGND _05262_ sg13g2_a21oi_1
X_11815_ _05250_ _05262_ VPWR VGND _05263_ sg13g2_nand2_1
X_11816_ _01056_ _05262_ _05263_ VPWR VGND _00742_ sg13g2_o21ai_1
X_11817_ _00785_ _00786_ _00007_ VPWR VGND _05264_ sg13g2_nand3_1
X_11818_ _05239_ _05264_ _05247_ VPWR VGND _05265_ sg13g2_a21oi_1
X_11819_ \atbs_core_0.uart_0.uart_rx_0.n2919_o\ _05250_ _05265_ VPWR VGND _00743_ sg13g2_mux2_1
X_11820_ _00788_ _05239_ _05247_ VPWR VGND _05266_ sg13g2_a21oi_1
X_11821_ \atbs_core_0.uart_0.uart_rx_0.n2921_o\ _05250_ _05266_ VPWR VGND _00744_ sg13g2_mux2_1
X_11822_ _00975_ _00815_ VPWR VGND _05267_ sg13g2_xor2_1
X_11823_ _01040_ _05267_ VPWR VGND _00745_ sg13g2_nor2_1
X_11824_ _00814_ VPWR VGND _05268_ sg13g2_inv_1
X_11825_ _00975_ _05268_ VPWR VGND _05269_ sg13g2_nand2_1
X_11826_ _00974_ _05269_ VPWR VGND _05270_ sg13g2_xnor2_1
X_11827_ _00978_ _05270_ VPWR VGND _00746_ sg13g2_and2_1
X_11828_ _00976_ _00815_ VPWR VGND _05271_ sg13g2_nand2_1
X_11829_ _00974_ _00975_ VPWR VGND _05272_ sg13g2_nand2_1
X_11830_ _00060_ _05272_ VPWR VGND _05273_ sg13g2_xor2_1
X_11831_ _05268_ _05273_ VPWR VGND _05274_ sg13g2_nand2_1
X_11832_ _05271_ _05274_ _01040_ VPWR VGND _00747_ sg13g2_a21oi_1
X_11833_ _02108_ VPWR VGND _05275_ sg13g2_buf_1
X_11834_ _01970_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ _05275_ VPWR VGND _00161_ sg13g2_mux2_1
X_11835_ _01902_ VPWR VGND _05276_ sg13g2_buf_1
X_11836_ _05276_ VPWR VGND _05277_ sg13g2_buf_1
X_11837_ _01928_ _05277_ VPWR VGND _05278_ sg13g2_nand2_1
X_11838_ _04156_ _02109_ _05278_ VPWR VGND _00162_ sg13g2_o21ai_1
X_11839_ _04124_ _02448_ VPWR VGND _05279_ sg13g2_nand2_1
X_11840_ _01936_ _04319_ _05279_ VPWR VGND _00163_ sg13g2_o21ai_1
X_11841_ _01914_ _05277_ VPWR VGND _05280_ sg13g2_nand2_1
X_11842_ _04142_ _02109_ _05280_ VPWR VGND _00164_ sg13g2_o21ai_1
X_11843_ _04148_ _02448_ VPWR VGND _05281_ sg13g2_nand2_1
X_11844_ _01911_ _04319_ _05281_ VPWR VGND _00165_ sg13g2_o21ai_1
X_11845_ _02447_ VPWR VGND _05282_ sg13g2_buf_1
X_11846_ _01905_ _04173_ _05282_ VPWR VGND _00166_ sg13g2_mux2_1
X_11847_ _04178_ _02448_ VPWR VGND _05283_ sg13g2_nand2_1
X_11848_ _02070_ _04319_ _05283_ VPWR VGND _00167_ sg13g2_o21ai_1
X_11849_ _02063_ _04123_ _05282_ VPWR VGND _00168_ sg13g2_mux2_1
X_11850_ _02447_ VPWR VGND _05284_ sg13g2_buf_1
X_11851_ _02081_ _04122_ _05284_ VPWR VGND _00169_ sg13g2_mux2_1
X_11852_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ _05277_ VPWR VGND _05285_ sg13g2_nand2_1
X_11853_ _01969_ _02109_ _05285_ VPWR VGND _00170_ sg13g2_o21ai_1
X_11854_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ _02448_ VPWR VGND _05286_ sg13g2_nand2_1
X_11855_ _02216_ _04319_ _05286_ VPWR VGND _00171_ sg13g2_o21ai_1
X_11856_ _02103_ VPWR VGND _05287_ sg13g2_buf_1
X_11857_ _02447_ VPWR VGND _05288_ sg13g2_buf_1
X_11858_ _02250_ _05288_ VPWR VGND _05289_ sg13g2_nand2_1
X_11859_ _01602_ _05287_ _05289_ VPWR VGND _00172_ sg13g2_o21ai_1
X_11860_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _05275_ VPWR VGND _00173_ sg13g2_mux2_1
X_11861_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ _05275_ VPWR VGND _00174_ sg13g2_mux2_1
X_11862_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ _05275_ VPWR VGND _00175_ sg13g2_mux2_1
X_11863_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _02229_ _05275_ VPWR VGND _00176_ sg13g2_mux2_1
X_11864_ _01920_ _02124_ _05275_ VPWR VGND _00177_ sg13g2_mux2_1
X_11865_ _01919_ _02125_ _05275_ VPWR VGND _00178_ sg13g2_mux2_1
X_11866_ _01924_ _02123_ _05275_ VPWR VGND _00179_ sg13g2_mux2_1
X_11867_ _01917_ _05288_ VPWR VGND _05290_ sg13g2_nand2_1
X_11868_ _02131_ _05287_ _05290_ VPWR VGND _00180_ sg13g2_o21ai_1
X_11869_ _01928_ _02122_ _05275_ VPWR VGND _00181_ sg13g2_mux2_1
X_11870_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[11]\ _05288_ VPWR VGND _05291_ sg13g2_nand2_1
X_11871_ _02121_ _05287_ _05291_ VPWR VGND _00182_ sg13g2_o21ai_1
X_11872_ _05117_ _05288_ VPWR VGND _05292_ sg13g2_nand2_1
X_11873_ _01664_ _05287_ _05292_ VPWR VGND _00183_ sg13g2_o21ai_1
X_11874_ _01914_ _05288_ VPWR VGND _05293_ sg13g2_nand2_1
X_11875_ _02120_ _05287_ _05293_ VPWR VGND _00184_ sg13g2_o21ai_1
X_11876_ _01910_ _05288_ VPWR VGND _05294_ sg13g2_nand2_1
X_11877_ _02118_ _05287_ _05294_ VPWR VGND _00185_ sg13g2_o21ai_1
X_11878_ _01905_ _02115_ _05275_ VPWR VGND _00186_ sg13g2_mux2_1
X_11879_ _02043_ _05288_ VPWR VGND _05295_ sg13g2_nand2_1
X_11880_ _02279_ _05287_ _05295_ VPWR VGND _00187_ sg13g2_o21ai_1
X_11881_ _01902_ VPWR VGND _05296_ sg13g2_buf_1
X_11882_ _05296_ VPWR VGND _05297_ sg13g2_buf_1
X_11883_ _02063_ _02150_ _05297_ VPWR VGND _00188_ sg13g2_mux2_1
X_11884_ _02081_ _05288_ VPWR VGND _05298_ sg13g2_nand2_1
X_11885_ _02114_ _05287_ _05298_ VPWR VGND _00189_ sg13g2_o21ai_1
X_11886_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ _05297_ VPWR VGND _00190_ sg13g2_mux2_1
X_11887_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ _05277_ VPWR VGND _05299_ sg13g2_nand2_1
X_11888_ _02216_ _02109_ _05299_ VPWR VGND _00191_ sg13g2_o21ai_1
X_11889_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _05288_ VPWR VGND _05300_ sg13g2_nand2_1
X_11890_ _02383_ _05287_ _05300_ VPWR VGND _00192_ sg13g2_o21ai_1
X_11891_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ _05288_ VPWR VGND _05301_ sg13g2_nand2_1
X_11892_ _02380_ _05287_ _05301_ VPWR VGND _00193_ sg13g2_o21ai_1
X_11893_ _01635_ _05277_ VPWR VGND _05302_ sg13g2_nand2_1
X_11894_ _02572_ _02109_ _05302_ VPWR VGND _00194_ sg13g2_o21ai_1
X_11895_ _02103_ VPWR VGND _05303_ sg13g2_buf_1
X_11896_ _02447_ VPWR VGND _05304_ sg13g2_buf_1
X_11897_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ _05304_ VPWR VGND _05305_ sg13g2_nand2_1
X_11898_ _02381_ _05303_ _05305_ VPWR VGND _00195_ sg13g2_o21ai_1
X_11899_ _02229_ _02390_ _05297_ VPWR VGND _00196_ sg13g2_mux2_1
X_11900_ _02124_ _02309_ _05297_ VPWR VGND _00197_ sg13g2_mux2_1
X_11901_ _02125_ _02310_ _05297_ VPWR VGND _00198_ sg13g2_mux2_1
X_11902_ _02123_ _02308_ _05297_ VPWR VGND _00199_ sg13g2_mux2_1
X_11903_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[9]\ _05304_ VPWR VGND _05306_ sg13g2_nand2_1
X_11904_ _02317_ _05303_ _05306_ VPWR VGND _00200_ sg13g2_o21ai_1
X_11905_ _02122_ _02307_ _05297_ VPWR VGND _00201_ sg13g2_mux2_1
X_11906_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[11]\ _05304_ VPWR VGND _05307_ sg13g2_nand2_1
X_11907_ _02306_ _05303_ _05307_ VPWR VGND _00202_ sg13g2_o21ai_1
X_11908_ _02119_ _05304_ VPWR VGND _05308_ sg13g2_nand2_1
X_11909_ _02305_ _05303_ _05308_ VPWR VGND _00203_ sg13g2_o21ai_1
X_11910_ _02327_ _05277_ VPWR VGND _05309_ sg13g2_nand2_1
X_11911_ _02118_ _02109_ _05309_ VPWR VGND _00204_ sg13g2_o21ai_1
X_11912_ _01632_ _05277_ VPWR VGND _05310_ sg13g2_nand2_1
X_11913_ _05134_ _02109_ _05310_ VPWR VGND _00205_ sg13g2_o21ai_1
X_11914_ _02115_ _05304_ VPWR VGND _05311_ sg13g2_nand2_1
X_11915_ _02335_ _05303_ _05311_ VPWR VGND _00206_ sg13g2_o21ai_1
X_11916_ _02108_ VPWR VGND _05312_ sg13g2_buf_1
X_11917_ _02339_ _05277_ VPWR VGND _05313_ sg13g2_nand2_1
X_11918_ _02279_ _05312_ _05313_ VPWR VGND _00207_ sg13g2_o21ai_1
X_11919_ _02150_ _02344_ _05297_ VPWR VGND _00208_ sg13g2_mux2_1
X_11920_ _02348_ _05277_ VPWR VGND _05314_ sg13g2_nand2_1
X_11921_ _02114_ _05312_ _05314_ VPWR VGND _00209_ sg13g2_o21ai_1
X_11922_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ _05297_ VPWR VGND _00210_ sg13g2_mux2_1
X_11923_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _05297_ VPWR VGND _00211_ sg13g2_mux2_1
X_11924_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ _05304_ VPWR VGND _05315_ sg13g2_nand2_1
X_11925_ _02539_ _05303_ _05315_ VPWR VGND _00212_ sg13g2_o21ai_1
X_11926_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ _05304_ VPWR VGND _05316_ sg13g2_nand2_1
X_11927_ _02538_ _05303_ _05316_ VPWR VGND _00213_ sg13g2_o21ai_1
X_11928_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ _05277_ VPWR VGND _05317_ sg13g2_nand2_1
X_11929_ _02381_ _05312_ _05317_ VPWR VGND _00214_ sg13g2_o21ai_1
X_11930_ _05296_ VPWR VGND _05318_ sg13g2_buf_1
X_11931_ _02390_ _02528_ _05318_ VPWR VGND _00215_ sg13g2_mux2_1
X_11932_ _01598_ VPWR VGND _05319_ sg13g2_inv_1
X_11933_ _02049_ _05304_ VPWR VGND _05320_ sg13g2_nand2_1
X_11934_ _05319_ _05303_ _05320_ VPWR VGND _00216_ sg13g2_o21ai_1
X_11935_ _02309_ _02461_ _05318_ VPWR VGND _00217_ sg13g2_mux2_1
X_11936_ _02310_ _02462_ _05318_ VPWR VGND _00218_ sg13g2_mux2_1
X_11937_ _02308_ _02466_ _05318_ VPWR VGND _00219_ sg13g2_mux2_1
X_11938_ _02460_ VPWR VGND _05321_ sg13g2_inv_1
X_11939_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[9]\ _05304_ VPWR VGND _05322_ sg13g2_nand2_1
X_11940_ _05321_ _05303_ _05322_ VPWR VGND _00220_ sg13g2_o21ai_1
X_11941_ _02307_ _02471_ _05318_ VPWR VGND _00221_ sg13g2_mux2_1
X_11942_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[11]\ _05304_ VPWR VGND _05323_ sg13g2_nand2_1
X_11943_ _02459_ _05303_ _05323_ VPWR VGND _00222_ sg13g2_o21ai_1
X_11944_ _05276_ VPWR VGND _05324_ sg13g2_buf_1
X_11945_ _02458_ _05324_ VPWR VGND _05325_ sg13g2_nand2_1
X_11946_ _02305_ _05312_ _05325_ VPWR VGND _00223_ sg13g2_o21ai_1
X_11947_ _02327_ _02457_ _05318_ VPWR VGND _00224_ sg13g2_mux2_1
X_11948_ _02103_ VPWR VGND _05326_ sg13g2_buf_1
X_11949_ _02447_ VPWR VGND _05327_ sg13g2_buf_1
X_11950_ _02328_ _05327_ VPWR VGND _05328_ sg13g2_nand2_1
X_11951_ _02484_ _05326_ _05328_ VPWR VGND _00225_ sg13g2_o21ai_1
X_11952_ _02339_ _05327_ VPWR VGND _05329_ sg13g2_nand2_1
X_11953_ _02455_ _05326_ _05329_ VPWR VGND _00226_ sg13g2_o21ai_1
X_11954_ _01596_ _05147_ _05284_ VPWR VGND _00227_ sg13g2_mux2_1
X_11955_ _02344_ _05327_ VPWR VGND _05330_ sg13g2_nand2_1
X_11956_ _02454_ _05326_ _05330_ VPWR VGND _00228_ sg13g2_o21ai_1
X_11957_ _02348_ _02453_ _05318_ VPWR VGND _00229_ sg13g2_mux2_1
X_11958_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ _05318_ VPWR VGND _00230_ sg13g2_mux2_1
X_11959_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _05327_ VPWR VGND _05331_ sg13g2_nand2_1
X_11960_ _02701_ _05326_ _05331_ VPWR VGND _00231_ sg13g2_o21ai_1
X_11961_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _05324_ VPWR VGND _05332_ sg13g2_nand2_1
X_11962_ _02539_ _05312_ _05332_ VPWR VGND _00232_ sg13g2_o21ai_1
X_11963_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _05324_ VPWR VGND _05333_ sg13g2_nand2_1
X_11964_ _02538_ _05312_ _05333_ VPWR VGND _00233_ sg13g2_o21ai_1
X_11965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ _05318_ VPWR VGND _00234_ sg13g2_mux2_1
X_11966_ _02528_ _02696_ _05318_ VPWR VGND _00235_ sg13g2_mux2_1
X_11967_ _05296_ VPWR VGND _05334_ sg13g2_buf_1
X_11968_ _02461_ _02612_ _05334_ VPWR VGND _00236_ sg13g2_mux2_1
X_11969_ _02462_ _02613_ _05334_ VPWR VGND _00237_ sg13g2_mux2_1
X_11970_ _01593_ _05324_ VPWR VGND _05335_ sg13g2_nand2_1
X_11971_ _03396_ _05312_ _05335_ VPWR VGND _00238_ sg13g2_o21ai_1
X_11972_ _02466_ _02611_ _05334_ VPWR VGND _00239_ sg13g2_mux2_1
X_11973_ _02460_ _05327_ VPWR VGND _05336_ sg13g2_nand2_1
X_11974_ _02610_ _05326_ _05336_ VPWR VGND _00240_ sg13g2_o21ai_1
X_11975_ _02471_ _02609_ _05334_ VPWR VGND _00241_ sg13g2_mux2_1
X_11976_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[11]\ _05327_ VPWR VGND _05337_ sg13g2_nand2_1
X_11977_ _02607_ _05326_ _05337_ VPWR VGND _00242_ sg13g2_o21ai_1
X_11978_ _02458_ _02605_ _05334_ VPWR VGND _00243_ sg13g2_mux2_1
X_11979_ _02457_ _02604_ _05334_ VPWR VGND _00244_ sg13g2_mux2_1
X_11980_ _02483_ _05327_ VPWR VGND _05338_ sg13g2_nand2_1
X_11981_ _02668_ _05326_ _05338_ VPWR VGND _00245_ sg13g2_o21ai_1
X_11982_ _02598_ _05324_ VPWR VGND _05339_ sg13g2_nand2_1
X_11983_ _02455_ _05312_ _05339_ VPWR VGND _00246_ sg13g2_o21ai_1
X_11984_ _02599_ _05324_ VPWR VGND _05340_ sg13g2_nand2_1
X_11985_ _02454_ _05312_ _05340_ VPWR VGND _00247_ sg13g2_o21ai_1
X_11986_ _02453_ _02641_ _05334_ VPWR VGND _00248_ sg13g2_mux2_1
X_11987_ _02086_ _05327_ VPWR VGND _05341_ sg13g2_nand2_1
X_11988_ _01694_ _05326_ _05341_ VPWR VGND _00249_ sg13g2_o21ai_1
X_11989_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ _05334_ VPWR VGND _00250_ sg13g2_mux2_1
X_11990_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[172]\ _05327_ VPWR VGND _05342_ sg13g2_nand2_1
X_11991_ _02848_ _05326_ _05342_ VPWR VGND _00251_ sg13g2_o21ai_1
X_11992_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _05327_ VPWR VGND _05343_ sg13g2_nand2_1
X_11993_ _02847_ _05326_ _05343_ VPWR VGND _00252_ sg13g2_o21ai_1
X_11994_ _02103_ VPWR VGND _05344_ sg13g2_buf_1
X_11995_ _02447_ VPWR VGND _05345_ sg13g2_buf_1
X_11996_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _05345_ VPWR VGND _05346_ sg13g2_nand2_1
X_11997_ _02846_ _05344_ _05346_ VPWR VGND _00253_ sg13g2_o21ai_1
X_11998_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ _05334_ VPWR VGND _00254_ sg13g2_mux2_1
X_11999_ _02696_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ _05334_ VPWR VGND _00255_ sg13g2_mux2_1
X_12000_ _05296_ VPWR VGND _05347_ sg13g2_buf_1
X_12001_ _02612_ _02789_ _05347_ VPWR VGND _00256_ sg13g2_mux2_1
X_12002_ _02613_ _02790_ _05347_ VPWR VGND _00257_ sg13g2_mux2_1
X_12003_ _02611_ _02788_ _05347_ VPWR VGND _00258_ sg13g2_mux2_1
X_12004_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[9]\ _05345_ VPWR VGND _05348_ sg13g2_nand2_1
X_12005_ _02798_ _05344_ _05348_ VPWR VGND _00259_ sg13g2_o21ai_1
X_12006_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ _05347_ VPWR VGND _00260_ sg13g2_mux2_1
X_12007_ _02609_ _02787_ _05347_ VPWR VGND _00261_ sg13g2_mux2_1
X_12008_ _02606_ _05345_ VPWR VGND _05349_ sg13g2_nand2_1
X_12009_ _02786_ _05344_ _05349_ VPWR VGND _00262_ sg13g2_o21ai_1
X_12010_ _02605_ _05345_ VPWR VGND _05350_ sg13g2_nand2_1
X_12011_ _02824_ _05344_ _05350_ VPWR VGND _00263_ sg13g2_o21ai_1
X_12012_ _02604_ _02808_ _05347_ VPWR VGND _00264_ sg13g2_mux2_1
X_12013_ _02603_ _05345_ VPWR VGND _05351_ sg13g2_nand2_1
X_12014_ _02780_ _05344_ _05351_ VPWR VGND _00265_ sg13g2_o21ai_1
X_12015_ _02598_ _02781_ _05347_ VPWR VGND _00266_ sg13g2_mux2_1
X_12016_ _02599_ _05345_ VPWR VGND _05352_ sg13g2_nand2_1
X_12017_ _02817_ _05344_ _05352_ VPWR VGND _00267_ sg13g2_o21ai_1
X_12018_ _02641_ _05345_ VPWR VGND _05353_ sg13g2_nand2_1
X_12019_ _02778_ _05344_ _05353_ VPWR VGND _00268_ sg13g2_o21ai_1
X_12020_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ _05347_ VPWR VGND _00269_ sg13g2_mux2_1
X_12021_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _05324_ VPWR VGND _05354_ sg13g2_nand2_1
X_12022_ _02848_ _05312_ _05354_ VPWR VGND _00270_ sg13g2_o21ai_1
X_12023_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _05345_ VPWR VGND _05355_ sg13g2_nand2_1
X_12024_ _03696_ _05344_ _05355_ VPWR VGND _00271_ sg13g2_o21ai_1
X_12025_ _02108_ VPWR VGND _05356_ sg13g2_buf_1
X_12026_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _05324_ VPWR VGND _05357_ sg13g2_nand2_1
X_12027_ _01797_ _05356_ _05357_ VPWR VGND _00272_ sg13g2_o21ai_1
X_12028_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ _05345_ VPWR VGND _05358_ sg13g2_nand2_1
X_12029_ _03040_ _05344_ _05358_ VPWR VGND _00273_ sg13g2_o21ai_1
X_12030_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _05324_ VPWR VGND _05359_ sg13g2_nand2_1
X_12031_ _02846_ _05356_ _05359_ VPWR VGND _00274_ sg13g2_o21ai_1
X_12032_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ _05347_ VPWR VGND _00275_ sg13g2_mux2_1
X_12033_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ _03030_ _05347_ VPWR VGND _00276_ sg13g2_mux2_1
X_12034_ _05296_ VPWR VGND _05360_ sg13g2_buf_1
X_12035_ _02789_ _02939_ _05360_ VPWR VGND _00277_ sg13g2_mux2_1
X_12036_ _02790_ _02940_ _05360_ VPWR VGND _00278_ sg13g2_mux2_1
X_12037_ _02788_ _02938_ _05360_ VPWR VGND _00279_ sg13g2_mux2_1
X_12038_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[9]\ _05345_ VPWR VGND _05361_ sg13g2_nand2_1
X_12039_ _02937_ _05344_ _05361_ VPWR VGND _00280_ sg13g2_o21ai_1
X_12040_ _02787_ _02935_ _05360_ VPWR VGND _00281_ sg13g2_mux2_1
X_12041_ _01107_ VPWR VGND _05362_ sg13g2_buf_1
X_12042_ _02589_ VPWR VGND _05363_ sg13g2_buf_1
X_12043_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[11]\ _05363_ VPWR VGND _05364_ sg13g2_nand2_1
X_12044_ _02934_ _05362_ _05364_ VPWR VGND _00282_ sg13g2_o21ai_1
X_12045_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[2]\ _05363_ VPWR VGND _05365_ sg13g2_nand2_1
X_12046_ _03695_ _05362_ _05365_ VPWR VGND _00283_ sg13g2_o21ai_1
X_12047_ _02954_ _05324_ VPWR VGND _05366_ sg13g2_nand2_1
X_12048_ _02824_ _05356_ _05366_ VPWR VGND _00284_ sg13g2_o21ai_1
X_12049_ _02808_ _02955_ _05360_ VPWR VGND _00285_ sg13g2_mux2_1
X_12050_ _02779_ _05363_ VPWR VGND _05367_ sg13g2_nand2_1
X_12051_ _02967_ _05362_ _05367_ VPWR VGND _00286_ sg13g2_o21ai_1
X_12052_ _02781_ _02930_ _05360_ VPWR VGND _00287_ sg13g2_mux2_1
X_12053_ _05276_ VPWR VGND _05368_ sg13g2_buf_1
X_12054_ _02929_ _05368_ VPWR VGND _05369_ sg13g2_nand2_1
X_12055_ _02817_ _05356_ _05369_ VPWR VGND _00288_ sg13g2_o21ai_1
X_12056_ _02928_ _05368_ VPWR VGND _05370_ sg13g2_nand2_1
X_12057_ _02778_ _05356_ _05370_ VPWR VGND _00289_ sg13g2_o21ai_1
X_12058_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ _05360_ VPWR VGND _00290_ sg13g2_mux2_1
X_12059_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _05363_ VPWR VGND _05371_ sg13g2_nand2_1
X_12060_ _03120_ _05362_ _05371_ VPWR VGND _00291_ sg13g2_o21ai_1
X_12061_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ _05363_ VPWR VGND _05372_ sg13g2_nand2_1
X_12062_ _03119_ _05362_ _05372_ VPWR VGND _00292_ sg13g2_o21ai_1
X_12063_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _05363_ VPWR VGND _05373_ sg13g2_nand2_1
X_12064_ _03118_ _05362_ _05373_ VPWR VGND _00293_ sg13g2_o21ai_1
X_12065_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _05363_ VPWR VGND _05374_ sg13g2_nand2_1
X_12066_ _03694_ _05362_ _05374_ VPWR VGND _00294_ sg13g2_o21ai_1
X_12067_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ _05360_ VPWR VGND _00295_ sg13g2_mux2_1
X_12068_ _03030_ _05363_ VPWR VGND _05375_ sg13g2_nand2_1
X_12069_ _03117_ _05362_ _05375_ VPWR VGND _00296_ sg13g2_o21ai_1
X_12070_ _02939_ _03098_ _05360_ VPWR VGND _00297_ sg13g2_mux2_1
X_12071_ _02940_ _03099_ _05360_ VPWR VGND _00298_ sg13g2_mux2_1
X_12072_ _05296_ VPWR VGND _05376_ sg13g2_buf_1
X_12073_ _02938_ _03103_ _05376_ VPWR VGND _00299_ sg13g2_mux2_1
X_12074_ _02936_ _05363_ VPWR VGND _05377_ sg13g2_nand2_1
X_12075_ _03148_ _05362_ _05377_ VPWR VGND _00300_ sg13g2_o21ai_1
X_12076_ _02935_ _03153_ _05376_ VPWR VGND _00301_ sg13g2_mux2_1
X_12077_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[11]\ _05363_ VPWR VGND _05378_ sg13g2_nand2_1
X_12078_ _03172_ _05362_ _05378_ VPWR VGND _00302_ sg13g2_o21ai_1
X_12079_ _02954_ _03171_ _05376_ VPWR VGND _00303_ sg13g2_mux2_1
X_12080_ _01107_ VPWR VGND _05379_ sg13g2_buf_1
X_12081_ _02589_ VPWR VGND _05380_ sg13g2_buf_1
X_12082_ _02955_ _05380_ VPWR VGND _05381_ sg13g2_nand2_1
X_12083_ _03202_ _05379_ _05381_ VPWR VGND _00304_ sg13g2_o21ai_1
X_12084_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ _05368_ VPWR VGND _05382_ sg13g2_nand2_1
X_12085_ _01785_ _05356_ _05382_ VPWR VGND _00305_ sg13g2_o21ai_1
X_12086_ _03194_ _05368_ VPWR VGND _05383_ sg13g2_nand2_1
X_12087_ _02967_ _05356_ _05383_ VPWR VGND _00306_ sg13g2_o21ai_1
X_12088_ _02930_ _03191_ _05376_ VPWR VGND _00307_ sg13g2_mux2_1
X_12089_ _02929_ _03219_ _05376_ VPWR VGND _00308_ sg13g2_mux2_1
X_12090_ _02928_ _03243_ _05376_ VPWR VGND _00309_ sg13g2_mux2_1
X_12091_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ _05376_ VPWR VGND _00310_ sg13g2_mux2_1
X_12092_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[229]\ _05380_ VPWR VGND _05384_ sg13g2_nand2_1
X_12093_ _03339_ _05379_ _05384_ VPWR VGND _00311_ sg13g2_o21ai_1
X_12094_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ _05380_ VPWR VGND _05385_ sg13g2_nand2_1
X_12095_ _03338_ _05379_ _05385_ VPWR VGND _00312_ sg13g2_o21ai_1
X_12096_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ _05380_ VPWR VGND _05386_ sg13g2_nand2_1
X_12097_ _03337_ _05379_ _05386_ VPWR VGND _00313_ sg13g2_o21ai_1
X_12098_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ _05376_ VPWR VGND _00314_ sg13g2_mux2_1
X_12099_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[233]\ _05380_ VPWR VGND _05387_ sg13g2_nand2_1
X_12100_ _03336_ _05379_ _05387_ VPWR VGND _00315_ sg13g2_o21ai_1
X_12101_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ _05380_ VPWR VGND _05388_ sg13g2_nand2_1
X_12102_ _03693_ _05379_ _05388_ VPWR VGND _00316_ sg13g2_o21ai_1
X_12103_ _03098_ _03280_ _05376_ VPWR VGND _00317_ sg13g2_mux2_1
X_12104_ _03099_ _03281_ _05376_ VPWR VGND _00318_ sg13g2_mux2_1
X_12105_ _05296_ VPWR VGND _05389_ sg13g2_buf_1
X_12106_ _03103_ _03279_ _05389_ VPWR VGND _00319_ sg13g2_mux2_1
X_12107_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[9]\ _05380_ VPWR VGND _05390_ sg13g2_nand2_1
X_12108_ _03278_ _05379_ _05390_ VPWR VGND _00320_ sg13g2_o21ai_1
X_12109_ _03153_ _03277_ _05389_ VPWR VGND _00321_ sg13g2_mux2_1
X_12110_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[11]\ _05380_ VPWR VGND _05391_ sg13g2_nand2_1
X_12111_ _03271_ _05379_ _05391_ VPWR VGND _00322_ sg13g2_o21ai_1
X_12112_ _03171_ _03270_ _05389_ VPWR VGND _00323_ sg13g2_mux2_1
X_12113_ _03272_ _05368_ VPWR VGND _05392_ sg13g2_nand2_1
X_12114_ _03202_ _05356_ _05392_ VPWR VGND _00324_ sg13g2_o21ai_1
X_12115_ _03194_ _03269_ _05389_ VPWR VGND _00325_ sg13g2_mux2_1
X_12116_ _03268_ VPWR VGND _05393_ sg13g2_inv_1
X_12117_ _03191_ _05380_ VPWR VGND _05394_ sg13g2_nand2_1
X_12118_ _05393_ _05379_ _05394_ VPWR VGND _00326_ sg13g2_o21ai_1
X_12119_ _01770_ _03616_ _05389_ VPWR VGND _00327_ sg13g2_mux2_1
X_12120_ _03219_ _03267_ _05389_ VPWR VGND _00328_ sg13g2_mux2_1
X_12121_ _03243_ _03306_ _05389_ VPWR VGND _00329_ sg13g2_mux2_1
X_12122_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ _05389_ VPWR VGND _00330_ sg13g2_mux2_1
X_12123_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[248]\ _05380_ VPWR VGND _05395_ sg13g2_nand2_1
X_12124_ _03467_ _05379_ _05395_ VPWR VGND _00331_ sg13g2_o21ai_1
X_12125_ _01107_ VPWR VGND _05396_ sg13g2_buf_1
X_12126_ _02589_ VPWR VGND _05397_ sg13g2_buf_1
X_12127_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ _05397_ VPWR VGND _05398_ sg13g2_nand2_1
X_12128_ _03466_ _05396_ _05398_ VPWR VGND _00332_ sg13g2_o21ai_1
X_12129_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ _05397_ VPWR VGND _05399_ sg13g2_nand2_1
X_12130_ _03465_ _05396_ _05399_ VPWR VGND _00333_ sg13g2_o21ai_1
X_12131_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _05389_ VPWR VGND _00334_ sg13g2_mux2_1
X_12132_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _05368_ VPWR VGND _05400_ sg13g2_nand2_1
X_12133_ _03336_ _05356_ _05400_ VPWR VGND _00335_ sg13g2_o21ai_1
X_12134_ _03280_ _03424_ _05389_ VPWR VGND _00336_ sg13g2_mux2_1
X_12135_ _05276_ VPWR VGND _05401_ sg13g2_buf_1
X_12136_ _03281_ _03425_ _05401_ VPWR VGND _00337_ sg13g2_mux2_1
X_12137_ _01762_ _03617_ _05401_ VPWR VGND _00338_ sg13g2_mux2_1
X_12138_ _03279_ _03423_ _05401_ VPWR VGND _00339_ sg13g2_mux2_1
X_12139_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[9]\ _05397_ VPWR VGND _05402_ sg13g2_nand2_1
X_12140_ _03422_ _05396_ _05402_ VPWR VGND _00340_ sg13g2_o21ai_1
X_12141_ _03277_ _03421_ _05401_ VPWR VGND _00341_ sg13g2_mux2_1
X_12142_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[11]\ _05397_ VPWR VGND _05403_ sg13g2_nand2_1
X_12143_ _03420_ _05396_ _05403_ VPWR VGND _00342_ sg13g2_o21ai_1
X_12144_ _03270_ _03419_ _05401_ VPWR VGND _00343_ sg13g2_mux2_1
X_12145_ _03272_ _03443_ _05401_ VPWR VGND _00344_ sg13g2_mux2_1
X_12146_ _03269_ _05397_ VPWR VGND _05404_ sg13g2_nand2_1
X_12147_ _03572_ _05396_ _05404_ VPWR VGND _00345_ sg13g2_o21ai_1
X_12148_ _03533_ _05368_ VPWR VGND _05405_ sg13g2_nand2_1
X_12149_ _05393_ _05356_ _05405_ VPWR VGND _00346_ sg13g2_o21ai_1
X_12150_ _03267_ _05397_ VPWR VGND _05406_ sg13g2_nand2_1
X_12151_ _03570_ _05396_ _05406_ VPWR VGND _00347_ sg13g2_o21ai_1
X_12152_ _03306_ _03555_ _05401_ VPWR VGND _00348_ sg13g2_mux2_1
X_12153_ _01607_ _03614_ _05401_ VPWR VGND _00349_ sg13g2_mux2_1
X_12154_ _01621_ _05397_ VPWR VGND _05407_ sg13g2_nand2_1
X_12155_ _03622_ _05396_ _05407_ VPWR VGND _00350_ sg13g2_o21ai_1
X_12156_ _02108_ VPWR VGND _05408_ sg13g2_buf_1
X_12157_ _03613_ _05368_ VPWR VGND _05409_ sg13g2_nand2_1
X_12158_ _01602_ _05408_ _05409_ VPWR VGND _00351_ sg13g2_o21ai_1
X_12159_ _01633_ _05397_ VPWR VGND _05410_ sg13g2_nand2_1
X_12160_ _03639_ _05396_ _05410_ VPWR VGND _00352_ sg13g2_o21ai_1
X_12161_ _02382_ _05397_ VPWR VGND _05411_ sg13g2_nand2_1
X_12162_ _01789_ _05396_ _05411_ VPWR VGND _00353_ sg13g2_o21ai_1
X_12163_ _01635_ _05397_ VPWR VGND _05412_ sg13g2_nand2_1
X_12164_ _03612_ _05396_ _05412_ VPWR VGND _00354_ sg13g2_o21ai_1
X_12165_ _01107_ VPWR VGND _05413_ sg13g2_buf_1
X_12166_ _02589_ VPWR VGND _05414_ sg13g2_buf_1
X_12167_ _01632_ _05414_ VPWR VGND _05415_ sg13g2_nand2_1
X_12168_ _03647_ _05413_ _05415_ VPWR VGND _00355_ sg13g2_o21ai_1
X_12169_ _03609_ _05368_ VPWR VGND _05416_ sg13g2_nand2_1
X_12170_ _05319_ _05408_ _05416_ VPWR VGND _00356_ sg13g2_o21ai_1
X_12171_ _01596_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[15]\ _05401_ VPWR VGND _00357_ sg13g2_mux2_1
X_12172_ _01593_ _03607_ _05401_ VPWR VGND _00358_ sg13g2_mux2_1
X_12173_ _03655_ _05368_ VPWR VGND _05417_ sg13g2_nand2_1
X_12174_ _01694_ _05408_ _05417_ VPWR VGND _00359_ sg13g2_o21ai_1
X_12175_ _05276_ VPWR VGND _05418_ sg13g2_buf_1
X_12176_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ _05418_ VPWR VGND _00360_ sg13g2_mux2_1
X_12177_ _05276_ VPWR VGND _05419_ sg13g2_buf_1
X_12178_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _05419_ VPWR VGND _05420_ sg13g2_nand2_1
X_12179_ _03696_ _05408_ _05420_ VPWR VGND _00361_ sg13g2_o21ai_1
X_12180_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ _05414_ VPWR VGND _05421_ sg13g2_nand2_1
X_12181_ _03862_ _05413_ _05421_ VPWR VGND _00362_ sg13g2_o21ai_1
X_12182_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _05419_ VPWR VGND _05422_ sg13g2_nand2_1
X_12183_ _03694_ _05408_ _05422_ VPWR VGND _00363_ sg13g2_o21ai_1
X_12184_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _05419_ VPWR VGND _05423_ sg13g2_nand2_1
X_12185_ _02222_ _05408_ _05423_ VPWR VGND _00364_ sg13g2_o21ai_1
X_12186_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ _05414_ VPWR VGND _05424_ sg13g2_nand2_1
X_12187_ _03861_ _05413_ _05424_ VPWR VGND _00365_ sg13g2_o21ai_1
X_12188_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[24]\ _05414_ VPWR VGND _05425_ sg13g2_nand2_1
X_12189_ _03860_ _05413_ _05425_ VPWR VGND _00366_ sg13g2_o21ai_1
X_12190_ _03616_ _03799_ _05418_ VPWR VGND _00367_ sg13g2_mux2_1
X_12191_ _03617_ _03800_ _05418_ VPWR VGND _00368_ sg13g2_mux2_1
X_12192_ _03614_ _03798_ _05418_ VPWR VGND _00369_ sg13g2_mux2_1
X_12193_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[9]\ _05414_ VPWR VGND _05426_ sg13g2_nand2_1
X_12194_ _03797_ _05413_ _05426_ VPWR VGND _00370_ sg13g2_o21ai_1
X_12195_ _03613_ _05414_ VPWR VGND _05427_ sg13g2_nand2_1
X_12196_ _03795_ _05413_ _05427_ VPWR VGND _00371_ sg13g2_o21ai_1
X_12197_ _03630_ _05414_ VPWR VGND _05428_ sg13g2_nand2_1
X_12198_ _03793_ _05413_ _05428_ VPWR VGND _00372_ sg13g2_o21ai_1
X_12199_ _03611_ _05414_ VPWR VGND _05429_ sg13g2_nand2_1
X_12200_ _03817_ _05413_ _05429_ VPWR VGND _00373_ sg13g2_o21ai_1
X_12201_ _03792_ _05419_ VPWR VGND _05430_ sg13g2_nand2_1
X_12202_ _03647_ _05408_ _05430_ VPWR VGND _00374_ sg13g2_o21ai_1
X_12203_ _01784_ _05414_ VPWR VGND _05431_ sg13g2_nand2_1
X_12204_ _01785_ _05413_ _05431_ VPWR VGND _00375_ sg13g2_o21ai_1
X_12205_ _03609_ _03819_ _05418_ VPWR VGND _00376_ sg13g2_mux2_1
X_12206_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[15]\ _05414_ VPWR VGND _05432_ sg13g2_nand2_1
X_12207_ _03826_ _05413_ _05432_ VPWR VGND _00377_ sg13g2_o21ai_1
X_12208_ _03607_ _03830_ _05418_ VPWR VGND _00378_ sg13g2_mux2_1
X_12209_ _01107_ VPWR VGND _05433_ sg13g2_buf_1
X_12210_ _02589_ VPWR VGND _05434_ sg13g2_buf_1
X_12211_ _03655_ _05434_ VPWR VGND _05435_ sg13g2_nand2_1
X_12212_ _03789_ _05433_ _05435_ VPWR VGND _00379_ sg13g2_o21ai_1
X_12213_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ _05418_ VPWR VGND _00380_ sg13g2_mux2_1
X_12214_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _05434_ VPWR VGND _05436_ sg13g2_nand2_1
X_12215_ _03995_ _05433_ _05436_ VPWR VGND _00381_ sg13g2_o21ai_1
X_12216_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[40]\ _05434_ VPWR VGND _05437_ sg13g2_nand2_1
X_12217_ _03994_ _05433_ _05437_ VPWR VGND _00382_ sg13g2_o21ai_1
X_12218_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _05434_ VPWR VGND _05438_ sg13g2_nand2_1
X_12219_ _03993_ _05433_ _05438_ VPWR VGND _00383_ sg13g2_o21ai_1
X_12220_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ _05419_ VPWR VGND _05439_ sg13g2_nand2_1
X_12221_ _03861_ _05408_ _05439_ VPWR VGND _00384_ sg13g2_o21ai_1
X_12222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[43]\ _05434_ VPWR VGND _05440_ sg13g2_nand2_1
X_12223_ _03992_ _05433_ _05440_ VPWR VGND _00385_ sg13g2_o21ai_1
X_12224_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ _05419_ VPWR VGND _05441_ sg13g2_nand2_1
X_12225_ _01980_ _05408_ _05441_ VPWR VGND _00386_ sg13g2_o21ai_1
X_12226_ _03799_ _03957_ _05418_ VPWR VGND _00387_ sg13g2_mux2_1
X_12227_ _03800_ _03958_ _05418_ VPWR VGND _00388_ sg13g2_mux2_1
X_12228_ _03798_ _03956_ _05418_ VPWR VGND _00389_ sg13g2_mux2_1
X_12229_ _03796_ _05434_ VPWR VGND _05442_ sg13g2_nand2_1
X_12230_ _03965_ _05433_ _05442_ VPWR VGND _00390_ sg13g2_o21ai_1
X_12231_ _03955_ _05419_ VPWR VGND _05443_ sg13g2_nand2_1
X_12232_ _03795_ _05408_ _05443_ VPWR VGND _00391_ sg13g2_o21ai_1
X_12233_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[11]\ _05434_ VPWR VGND _05444_ sg13g2_nand2_1
X_12234_ _03954_ _05433_ _05444_ VPWR VGND _00392_ sg13g2_o21ai_1
X_12235_ _03816_ _05434_ VPWR VGND _05445_ sg13g2_nand2_1
X_12236_ _03953_ _05433_ _05445_ VPWR VGND _00393_ sg13g2_o21ai_1
X_12237_ _05276_ VPWR VGND _05446_ sg13g2_buf_1
X_12238_ _03792_ _03978_ _05446_ VPWR VGND _00394_ sg13g2_mux2_1
X_12239_ _03819_ _05434_ VPWR VGND _05447_ sg13g2_nand2_1
X_12240_ _04059_ _05433_ _05447_ VPWR VGND _00395_ sg13g2_o21ai_1
X_12241_ _02108_ VPWR VGND _05448_ sg13g2_buf_1
X_12242_ _04062_ _05419_ VPWR VGND _05449_ sg13g2_nand2_1
X_12243_ _03826_ _05448_ _05449_ VPWR VGND _00396_ sg13g2_o21ai_1
X_12244_ _01770_ _05419_ VPWR VGND _05450_ sg13g2_nand2_1
X_12245_ _01983_ _05448_ _05450_ VPWR VGND _00397_ sg13g2_o21ai_1
X_12246_ _03830_ _04078_ _05446_ VPWR VGND _00398_ sg13g2_mux2_1
X_12247_ _03788_ _05434_ VPWR VGND _05451_ sg13g2_nand2_1
X_12248_ _04113_ _05433_ _05451_ VPWR VGND _00399_ sg13g2_o21ai_1
X_12249_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ _05446_ VPWR VGND _00400_ sg13g2_mux2_1
X_12250_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _05419_ VPWR VGND _05452_ sg13g2_nand2_1
X_12251_ _03995_ _05448_ _05452_ VPWR VGND _00401_ sg13g2_o21ai_1
X_12252_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ _02593_ VPWR VGND _05453_ sg13g2_nand2_1
X_12253_ _03994_ _05448_ _05453_ VPWR VGND _00402_ sg13g2_o21ai_1
X_12254_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _02593_ VPWR VGND _05454_ sg13g2_nand2_1
X_12255_ _03993_ _05448_ _05454_ VPWR VGND _00403_ sg13g2_o21ai_1
X_12256_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _05446_ VPWR VGND _00404_ sg13g2_mux2_1
X_12257_ _04211_ _02593_ VPWR VGND _05455_ sg13g2_nand2_1
X_12258_ _03992_ _05448_ _05455_ VPWR VGND _00405_ sg13g2_o21ai_1
X_12259_ _03957_ _04128_ _05446_ VPWR VGND _00406_ sg13g2_mux2_1
X_12260_ _03958_ _04129_ _05446_ VPWR VGND _00407_ sg13g2_mux2_1
X_12261_ _01762_ _02593_ VPWR VGND _05456_ sg13g2_nand2_1
X_12262_ _05194_ _05448_ _05456_ VPWR VGND _00408_ sg13g2_o21ai_1
X_12263_ _03956_ _04127_ _05446_ VPWR VGND _00409_ sg13g2_mux2_1
X_12264_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[9]\ _02590_ VPWR VGND _05457_ sg13g2_nand2_1
X_12265_ _04134_ _05282_ _05457_ VPWR VGND _00410_ sg13g2_o21ai_1
X_12266_ _03955_ _02590_ VPWR VGND _05458_ sg13g2_nand2_1
X_12267_ _04156_ _05282_ _05458_ VPWR VGND _00411_ sg13g2_o21ai_1
X_12268_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[11]\ _02590_ VPWR VGND _05459_ sg13g2_nand2_1
X_12269_ _04125_ _05282_ _05459_ VPWR VGND _00412_ sg13g2_o21ai_1
X_12270_ _03952_ _02590_ VPWR VGND _05460_ sg13g2_nand2_1
X_12271_ _04142_ _05282_ _05460_ VPWR VGND _00413_ sg13g2_o21ai_1
X_12272_ _03978_ _04148_ _05446_ VPWR VGND _00414_ sg13g2_mux2_1
X_12273_ _04173_ _02593_ VPWR VGND _05461_ sg13g2_nand2_1
X_12274_ _04059_ _05448_ _05461_ VPWR VGND _00415_ sg13g2_o21ai_1
X_12275_ _04062_ _04178_ _05446_ VPWR VGND _00416_ sg13g2_mux2_1
X_12276_ _04078_ _04123_ _05446_ VPWR VGND _00417_ sg13g2_mux2_1
X_12277_ _04122_ _02593_ VPWR VGND _05462_ sg13g2_nand2_1
X_12278_ _04113_ _05448_ _05462_ VPWR VGND _00418_ sg13g2_o21ai_1
X_12279_ _01607_ _02593_ VPWR VGND _05463_ sg13g2_nand2_1
X_12280_ _04239_ _05448_ _05463_ VPWR VGND _00419_ sg13g2_o21ai_1
X_12281_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ _02590_ VPWR VGND _05464_ sg13g2_nand2_1
X_12282_ _01969_ _05282_ _05464_ VPWR VGND _00420_ sg13g2_o21ai_1
X_12283_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _05284_ VPWR VGND _00421_ sg13g2_mux2_1
X_12284_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ _05284_ VPWR VGND _00422_ sg13g2_mux2_1
X_12285_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _05284_ VPWR VGND _00423_ sg13g2_mux2_1
X_12286_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _05284_ VPWR VGND _00424_ sg13g2_mux2_1
X_12287_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _04211_ _05284_ VPWR VGND _00425_ sg13g2_mux2_1
X_12288_ _01920_ _04128_ _05284_ VPWR VGND _00426_ sg13g2_mux2_1
X_12289_ _01919_ _04129_ _05284_ VPWR VGND _00427_ sg13g2_mux2_1
X_12290_ _01924_ _04127_ _05284_ VPWR VGND _00428_ sg13g2_mux2_1
X_12291_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[9]\ _02590_ VPWR VGND _05465_ sg13g2_nand2_1
X_12292_ _01918_ _05282_ _05465_ VPWR VGND _00429_ sg13g2_o21ai_1
X_12293_ _05100_ _02590_ VPWR VGND _05466_ sg13g2_nand2_1
X_12294_ _01622_ _05282_ _05466_ VPWR VGND _00430_ sg13g2_o21ai_1
X_12295_ \atbs_core_0.dac_control_0.n1495_o\ VPWR VGND _05467_ sg13g2_inv_1
X_12296_ \atbs_core_0.dac_control_0.dac_init_value[1]\ _05467_ VPWR VGND _05468_ sg13g2_nor2_1
X_12297_ _05467_ _04345_ _05468_ VPWR VGND _00476_ sg13g2_a21oi_1
X_12298_ \atbs_core_0.dac_control_0.n1495_o\ VPWR VGND _05469_ sg13g2_buf_1
X_12299_ _05469_ \atbs_core_0.dac_control_0.dac_init_value[2]\ VPWR VGND _05470_ sg13g2_nand2_1
X_12300_ _05469_ _04368_ _05470_ VPWR VGND _00477_ sg13g2_o21ai_1
X_12301_ _05469_ \atbs_core_0.dac_control_0.dac_init_value[3]\ VPWR VGND _05471_ sg13g2_nand2_1
X_12302_ _05469_ _04357_ _05471_ VPWR VGND _00478_ sg13g2_o21ai_1
X_12303_ _05469_ \atbs_core_0.dac_control_0.dac_init_value[4]\ VPWR VGND _05472_ sg13g2_nand2_1
X_12304_ _05469_ _04346_ _05472_ VPWR VGND _00479_ sg13g2_o21ai_1
X_12305_ \atbs_core_0.dac_control_0.dac_init_value[5]\ _04400_ _05467_ VPWR VGND _00480_ sg13g2_mux2_1
X_12306_ \atbs_core_0.dac_control_0.dac_init_value[6]\ _04406_ _05467_ VPWR VGND _00481_ sg13g2_mux2_1
X_12307_ \atbs_core_0.dac_control_0.dac_init_value[7]\ _05469_ VPWR VGND _00482_ sg13g2_nand2b_1
X_12308_ _05469_ \atbs_core_0.dac_control_0.dac_init_value[8]\ VPWR VGND _00483_ sg13g2_and2_1
X_12309_ \atbs_core_0.dac_control_1.dac_init_value[7]\ \atbs_core_0.dac_control_1.n1629_o\ VPWR VGND _00502_ sg13g2_nand2b_1
X_12310_ _00847_ _00848_ VPWR VGND _05473_ sg13g2_nor2_1
X_12311_ _00841_ _05473_ VPWR VGND _05474_ sg13g2_and2_1
X_12312_ _05474_ VPWR VGND _05475_ sg13g2_buf_1
X_12313_ _00846_ _05475_ VPWR VGND _05476_ sg13g2_nand2b_1
X_12314_ _01035_ _01070_ _01072_ _05476_ VPWR VGND 
+ _05477_
+ sg13g2_a22oi_1
X_12315_ _00027_ VPWR VGND _05478_ sg13g2_inv_1
X_12316_ _00842_ _05478_ VPWR VGND _05479_ sg13g2_nor2_1
X_12317_ _05477_ _05479_ VPWR VGND _05480_ sg13g2_nor2b_1
X_12318_ _00841_ _00851_ _01094_ VPWR VGND _05481_ sg13g2_a21oi_1
X_12319_ _01074_ _05481_ VPWR VGND _05482_ sg13g2_nand2b_1
X_12320_ _00843_ _05069_ _01092_ VPWR VGND _05483_ sg13g2_nor3_1
X_12321_ _00846_ _05475_ _00844_ VPWR VGND _05484_ sg13g2_a21oi_1
X_12322_ _05483_ _05484_ VPWR VGND _05485_ sg13g2_nor2_1
X_12323_ _01035_ _01072_ VPWR VGND _05486_ sg13g2_nand2_1
X_12324_ _01069_ _05485_ _05486_ VPWR VGND _05487_ sg13g2_o21ai_1
X_12325_ _04985_ _05487_ VPWR VGND _05488_ sg13g2_and2_1
X_12326_ _05480_ _05482_ _05488_ VPWR VGND _00121_ sg13g2_nor3_1
X_12327_ _05236_ VPWR VGND _05489_ sg13g2_inv_1
X_12328_ _00971_ uart_rx_i _05489_ _00956_ VPWR VGND 
+ _00123_
+ sg13g2_a22oi_1
X_12329_ _00817_ _00815_ VPWR VGND _05490_ sg13g2_nor2_1
X_12330_ _00819_ \atbs_core_0.uart_0.uart_tx_0.n2721_o\ _00031_ _05490_ VPWR VGND 
+ _00124_
+ sg13g2_a22oi_1
X_12331_ _01138_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1345_o\ sg13g2_inv_1
X_12332_ _00051_ _01134_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1348_o\ sg13g2_nor2_1
X_12333_ _02596_ VPWR VGND _05491_ sg13g2_inv_1
X_12334_ _00075_ VPWR VGND _05492_ sg13g2_buf_1
X_12335_ _05492_ VPWR VGND _05493_ sg13g2_inv_1
X_12336_ _02776_ VPWR VGND _05494_ sg13g2_inv_1
X_12337_ _00074_ VPWR VGND _05495_ sg13g2_buf_1
X_12338_ _03261_ VPWR VGND _05496_ sg13g2_inv_1
X_12339_ _00072_ VPWR VGND _05497_ sg13g2_buf_1
X_12340_ _05497_ VPWR VGND _05498_ sg13g2_inv_1
X_12341_ _03591_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2931_o\ VPWR VGND _05499_ sg13g2_nor2b_1
X_12342_ _05499_ VPWR VGND _05500_ sg13g2_buf_1
X_12343_ _03264_ _03415_ VPWR VGND _05501_ sg13g2_nor2b_1
X_12344_ _03263_ _05500_ _05501_ VPWR VGND _05502_ sg13g2_nand3_1
X_12345_ _03263_ _05498_ _05502_ VPWR VGND _05503_ sg13g2_o21ai_1
X_12346_ _00073_ VPWR VGND _05504_ sg13g2_buf_1
X_12347_ _05500_ _05504_ _03264_ VPWR VGND _05505_ sg13g2_mux2_1
X_12348_ _03591_ _05504_ VPWR VGND _05506_ sg13g2_nor2b_1
X_12349_ _05505_ _05506_ _03415_ VPWR VGND _05507_ sg13g2_mux2_1
X_12350_ _05507_ VPWR VGND _05508_ sg13g2_buf_1
X_12351_ _05496_ _05498_ VPWR VGND _05509_ sg13g2_nor2_1
X_12352_ _05496_ _05503_ _05508_ _05509_ VPWR VGND 
+ _05510_
+ sg13g2_a22oi_1
X_12353_ _00071_ VPWR VGND _05511_ sg13g2_buf_1
X_12354_ _03093_ _05511_ VPWR VGND _05512_ sg13g2_nand2_1
X_12355_ _03261_ _03263_ _05500_ _05501_ VPWR VGND 
+ _05513_
+ sg13g2_and4_1
X_12356_ _05513_ VPWR VGND _05514_ sg13g2_buf_1
X_12357_ _05511_ _05514_ _03090_ VPWR VGND _05515_ sg13g2_mux2_1
X_12358_ _03094_ _05515_ VPWR VGND _05516_ sg13g2_nand2_1
X_12359_ _05510_ _05512_ _05516_ VPWR VGND _05517_ sg13g2_o21ai_1
X_12360_ _05495_ _05517_ VPWR VGND _05518_ sg13g2_or2_1
X_12361_ _03090_ _05511_ _05514_ VPWR VGND _05519_ sg13g2_nor3_1
X_12362_ _05496_ _05503_ _05508_ _05509_ _03089_ VPWR 
+ VGND
+ _05520_ sg13g2_a221oi_1
X_12363_ _03093_ _05519_ _05520_ VPWR VGND _05521_ sg13g2_or3_1
X_12364_ _05500_ _05501_ _05497_ VPWR VGND _05522_ sg13g2_a21oi_1
X_12365_ _03097_ _05522_ VPWR VGND _05523_ sg13g2_and2_1
X_12366_ _03416_ _03591_ VPWR VGND _05524_ sg13g2_nor2_1
X_12367_ _03416_ _05505_ _05524_ _05504_ _03097_ VPWR 
+ VGND
+ _05525_ sg13g2_a221oi_1
X_12368_ _03261_ _05523_ _05525_ VPWR VGND _05526_ sg13g2_nor3_1
X_12369_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2931_o\ VPWR VGND _05527_ sg13g2_inv_1
X_12370_ _03415_ _03264_ VPWR VGND _05528_ sg13g2_or2_1
X_12371_ _05527_ _05528_ _03591_ VPWR VGND _05529_ sg13g2_a21oi_1
X_12372_ _05504_ _05528_ VPWR VGND _05530_ sg13g2_and2_1
X_12373_ _05529_ _05530_ VPWR VGND _05531_ sg13g2_nor2_1
X_12374_ _05496_ _05522_ _05531_ VPWR VGND _05532_ sg13g2_nor3_1
X_12375_ _05511_ _05514_ VPWR VGND _05533_ sg13g2_nor2_1
X_12376_ _03094_ _05533_ VPWR VGND _05534_ sg13g2_nor2_1
X_12377_ _05526_ _05532_ _05534_ VPWR VGND _05535_ sg13g2_o21ai_1
X_12378_ _05494_ _05521_ _05535_ VPWR VGND _05536_ sg13g2_nand3_1
X_12379_ _05494_ _05518_ _05536_ VPWR VGND _05537_ sg13g2_o21ai_1
X_12380_ _05511_ VPWR VGND _05538_ sg13g2_inv_1
X_12381_ _03089_ _05538_ _05510_ VPWR VGND _05539_ sg13g2_and3_1
X_12382_ _03089_ _05526_ _05532_ VPWR VGND _05540_ sg13g2_nor3_1
X_12383_ _03093_ _05539_ _05540_ VPWR VGND _05541_ sg13g2_nor3_1
X_12384_ _05538_ _05510_ VPWR VGND _05542_ sg13g2_nand2_1
X_12385_ _03416_ _05505_ _05524_ _05504_ _05497_ VPWR 
+ VGND
+ _05543_ sg13g2_a221oi_1
X_12386_ _03097_ _05529_ _05530_ VPWR VGND _05544_ sg13g2_nor3_1
X_12387_ _03097_ _05543_ _05544_ VPWR VGND _05545_ sg13g2_a21oi_1
X_12388_ _03264_ _03591_ VPWR VGND _05546_ sg13g2_and2_1
X_12389_ _05546_ VPWR VGND _05547_ sg13g2_buf_1
X_12390_ _05496_ _05547_ VPWR VGND _05548_ sg13g2_nor2_1
X_12391_ _05543_ _05548_ VPWR VGND _05549_ sg13g2_nor2b_1
X_12392_ _05496_ _05545_ _05549_ VPWR VGND _05550_ sg13g2_a21o_1
X_12393_ _03093_ _05542_ _05550_ VPWR VGND _05551_ sg13g2_and3_1
X_12394_ _05551_ VPWR VGND _05552_ sg13g2_buf_1
X_12395_ _05541_ _05552_ _05518_ VPWR VGND _05553_ sg13g2_o21ai_1
X_12396_ _05537_ _05553_ _02926_ VPWR VGND _05554_ sg13g2_mux2_1
X_12397_ _02926_ VPWR VGND _05555_ sg13g2_inv_1
X_12398_ _05555_ VPWR VGND _05556_ sg13g2_buf_1
X_12399_ _05495_ VPWR VGND _05557_ sg13g2_inv_1
X_12400_ _05541_ _05552_ VPWR VGND _05558_ sg13g2_nor2_1
X_12401_ _05497_ _05508_ VPWR VGND _05559_ sg13g2_or2_1
X_12402_ _05496_ _05545_ _05548_ _05559_ _05511_ VPWR 
+ VGND
+ _05560_ sg13g2_a221oi_1
X_12403_ _03261_ _03097_ VPWR VGND _05561_ sg13g2_nor2_1
X_12404_ _05497_ _05561_ VPWR VGND _05562_ sg13g2_nor2_1
X_12405_ _05547_ _05561_ _05562_ _05531_ VPWR VGND 
+ _05563_
+ sg13g2_a22oi_1
X_12406_ _05563_ VPWR VGND _05564_ sg13g2_buf_1
X_12407_ _03090_ _05564_ VPWR VGND _05565_ sg13g2_nand2_1
X_12408_ _03090_ _05560_ _05565_ VPWR VGND _05566_ sg13g2_o21ai_1
X_12409_ _05547_ _05562_ VPWR VGND _05567_ sg13g2_and2_1
X_12410_ _05567_ VPWR VGND _05568_ sg13g2_buf_1
X_12411_ _03094_ _05560_ _05568_ VPWR VGND _05569_ sg13g2_nor3_1
X_12412_ _03094_ _05566_ _05569_ VPWR VGND _05570_ sg13g2_a21oi_1
X_12413_ _05557_ _05558_ _05570_ VPWR VGND _05571_ sg13g2_a21oi_1
X_12414_ _05494_ _05495_ _05541_ _05552_ VPWR VGND 
+ _05572_
+ sg13g2_nor4_1
X_12415_ _03090_ _05511_ _05526_ _05532_ VPWR VGND 
+ _05573_
+ sg13g2_nor4_1
X_12416_ _05496_ _05545_ _05548_ _05559_ _03089_ VPWR 
+ VGND
+ _05574_ sg13g2_a221oi_1
X_12417_ _03093_ _05573_ _05574_ VPWR VGND _05575_ sg13g2_nor3_1
X_12418_ _05526_ _05532_ VPWR VGND _05576_ sg13g2_nor2_1
X_12419_ _03093_ _05564_ VPWR VGND _05577_ sg13g2_nand2_1
X_12420_ _05538_ _05576_ _05577_ VPWR VGND _05578_ sg13g2_a21oi_1
X_12421_ _02776_ _05575_ _05578_ VPWR VGND _05579_ sg13g2_nor3_1
X_12422_ _05572_ _05579_ _05556_ VPWR VGND _05580_ sg13g2_o21ai_1
X_12423_ _05556_ _05571_ _05580_ VPWR VGND _05581_ sg13g2_o21ai_1
X_12424_ _05493_ _05554_ _05581_ VPWR VGND _05582_ sg13g2_a21oi_1
X_12425_ _05556_ _05575_ _05578_ VPWR VGND _05583_ sg13g2_nor3_1
X_12426_ _05521_ _05535_ VPWR VGND _05584_ sg13g2_nand2_1
X_12427_ _05555_ _05494_ VPWR VGND _05585_ sg13g2_nand2_1
X_12428_ _05495_ _05584_ _05585_ VPWR VGND _05586_ sg13g2_o21ai_1
X_12429_ _02926_ _02776_ VPWR VGND _05587_ sg13g2_nor2_1
X_12430_ _05541_ _05552_ _05587_ VPWR VGND _05588_ sg13g2_o21ai_1
X_12431_ _05583_ _05586_ _05588_ VPWR VGND _05589_ sg13g2_o21ai_1
X_12432_ _02766_ _02759_ VPWR VGND _05590_ sg13g2_nor2_1
X_12433_ _05590_ VPWR VGND _05591_ sg13g2_buf_1
X_12434_ _02767_ _02759_ VPWR VGND _05592_ sg13g2_nand2_1
X_12435_ _05493_ _05554_ _05592_ VPWR VGND _05593_ sg13g2_a21oi_1
X_12436_ _05589_ _05591_ _05593_ VPWR VGND _05594_ sg13g2_a21o_1
X_12437_ _02766_ _05582_ _05594_ VPWR VGND _05595_ sg13g2_a21o_1
X_12438_ _00076_ VPWR VGND _05596_ sg13g2_inv_1
X_12439_ _05493_ _05554_ VPWR VGND _05597_ sg13g2_nor2_1
X_12440_ _05492_ _02759_ VPWR VGND _05598_ sg13g2_nor2b_1
X_12441_ _02776_ _05517_ VPWR VGND _05599_ sg13g2_nor2_1
X_12442_ _02776_ _05557_ _05599_ VPWR VGND _05600_ sg13g2_a21oi_1
X_12443_ _05556_ _05557_ VPWR VGND _05601_ sg13g2_nor2_1
X_12444_ _05556_ _05600_ _05601_ _05584_ _02759_ VPWR 
+ VGND
+ _05602_ sg13g2_a221oi_1
X_12445_ _02766_ _05598_ _05602_ VPWR VGND _05603_ sg13g2_nor3_1
X_12446_ _02766_ _05597_ _05603_ VPWR VGND _05604_ sg13g2_a21oi_1
X_12447_ _02596_ _02592_ VPWR VGND _05605_ sg13g2_nor2_1
X_12448_ _05596_ _05604_ _05605_ VPWR VGND _05606_ sg13g2_a21oi_1
X_12449_ _05491_ _05595_ _05606_ VPWR VGND _05607_ sg13g2_o21ai_1
X_12450_ _05556_ _05553_ VPWR VGND _05608_ sg13g2_or2_1
X_12451_ _02926_ _05537_ _05608_ VPWR VGND _05609_ sg13g2_o21ai_1
X_12452_ _05556_ _05600_ _05601_ _05584_ _05492_ VPWR 
+ VGND
+ _05610_ sg13g2_a221oi_1
X_12453_ _02767_ _05610_ VPWR VGND _05611_ sg13g2_nor2_1
X_12454_ _05592_ _05610_ VPWR VGND _05612_ sg13g2_nor2_1
X_12455_ _05609_ _05591_ _05611_ _05589_ _05612_ VPWR 
+ VGND
+ _05613_ sg13g2_a221oi_1
X_12456_ _05613_ VPWR VGND _05614_ sg13g2_buf_1
X_12457_ _05614_ _05605_ VPWR VGND _05615_ sg13g2_nand2b_1
X_12458_ _05607_ _05615_ VPWR VGND _05616_ sg13g2_and2_1
X_12459_ _05616_ VPWR VGND _05617_ sg13g2_buf_1
X_12460_ _02592_ _05604_ VPWR VGND _05618_ sg13g2_nor2b_1
X_12461_ _02592_ _05596_ _05618_ VPWR VGND _05619_ sg13g2_a21oi_1
X_12462_ _05491_ _05596_ _05614_ VPWR VGND _05620_ sg13g2_nor3_1
X_12463_ _05491_ _05619_ _05620_ VPWR VGND _05621_ sg13g2_a21oi_1
X_12464_ _05617_ _05621_ _02451_ VPWR VGND _05622_ sg13g2_mux2_1
X_12465_ _02302_ _05622_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[48]\ sg13g2_or2_1
X_12466_ _05492_ _05589_ VPWR VGND _05623_ sg13g2_nor2_1
X_12467_ _03093_ _03089_ VPWR VGND _05624_ sg13g2_nor2_1
X_12468_ _05511_ _05564_ _05624_ VPWR VGND _05625_ sg13g2_nor3_1
X_12469_ _05568_ _05624_ _05625_ VPWR VGND _05626_ sg13g2_a21o_1
X_12470_ _05556_ _05626_ VPWR VGND _05627_ sg13g2_or2_1
X_12471_ _05556_ _02776_ VPWR VGND _05628_ sg13g2_nand2_1
X_12472_ _05495_ _05575_ _05578_ VPWR VGND _05629_ sg13g2_nor3_1
X_12473_ _05627_ _05628_ _05629_ VPWR VGND _05630_ sg13g2_a21o_1
X_12474_ _05570_ _05585_ _05630_ VPWR VGND _05631_ sg13g2_o21ai_1
X_12475_ _05631_ VPWR VGND _05632_ sg13g2_buf_1
X_12476_ _05623_ _05632_ VPWR VGND _05633_ sg13g2_nand2b_1
X_12477_ _05581_ _05623_ _02759_ VPWR VGND _05634_ sg13g2_mux2_1
X_12478_ _05633_ _05634_ _02767_ VPWR VGND _05635_ sg13g2_mux2_1
X_12479_ _05596_ _05614_ _05491_ VPWR VGND _05636_ sg13g2_a21o_1
X_12480_ _05491_ _02592_ VPWR VGND _05637_ sg13g2_nand2_1
X_12481_ _05596_ _05614_ _05637_ VPWR VGND _05638_ sg13g2_a21oi_1
X_12482_ _05595_ _05605_ _05638_ VPWR VGND _05639_ sg13g2_a21oi_1
X_12483_ _05635_ _05636_ _05639_ VPWR VGND _05640_ sg13g2_o21ai_1
X_12484_ _05640_ VPWR VGND _05641_ sg13g2_buf_1
X_12485_ _02450_ _02302_ VPWR VGND _05642_ sg13g2_nor2_1
X_12486_ _02302_ _05621_ _05642_ _05617_ VPWR VGND 
+ _05643_
+ sg13g2_a22oi_1
X_12487_ _02451_ _05641_ _05643_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[49]\ sg13g2_o21ai_1
X_12488_ _05635_ VPWR VGND _05644_ sg13g2_inv_1
X_12489_ _02766_ _05582_ _05594_ VPWR VGND _05645_ sg13g2_a21oi_1
X_12490_ _05495_ _05587_ VPWR VGND _05646_ sg13g2_nor2_1
X_12491_ _05587_ _05626_ VPWR VGND _05647_ sg13g2_and2_1
X_12492_ _05570_ _05646_ _05647_ VPWR VGND _05648_ sg13g2_a21o_1
X_12493_ _05648_ VPWR VGND _05649_ sg13g2_buf_1
X_12494_ _02767_ _05649_ VPWR VGND _05650_ sg13g2_or2_1
X_12495_ _05493_ _05581_ _05592_ _05650_ VPWR VGND 
+ _05651_
+ sg13g2_a22oi_1
X_12496_ _05591_ _05632_ _05651_ VPWR VGND _05652_ sg13g2_a21oi_1
X_12497_ _05596_ _05645_ _05652_ VPWR VGND _05653_ sg13g2_a21oi_1
X_12498_ _05596_ _05645_ _05637_ VPWR VGND _05654_ sg13g2_a21oi_1
X_12499_ _05605_ _05644_ _05653_ _02596_ _05654_ VPWR 
+ VGND
+ _05655_ sg13g2_a221oi_1
X_12500_ _05655_ VPWR VGND _05656_ sg13g2_buf_1
X_12501_ _02451_ _02303_ VPWR VGND _05657_ sg13g2_nand2_1
X_12502_ _05657_ _05641_ VPWR VGND _05658_ sg13g2_nor2_1
X_12503_ _02302_ _05617_ _05656_ _02450_ _05658_ VPWR 
+ VGND
+ _05659_ sg13g2_a221oi_1
X_12504_ _05659_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[50]\ sg13g2_inv_1
X_12505_ _05492_ _05591_ _05632_ VPWR VGND _05660_ sg13g2_nor3_1
X_12506_ _05591_ _05649_ VPWR VGND _05661_ sg13g2_nand2_1
X_12507_ _05660_ _02596_ _05661_ VPWR VGND _05662_ sg13g2_nand3b_1
X_12508_ _05596_ _05635_ _05637_ _05662_ VPWR VGND 
+ _05663_
+ sg13g2_a22oi_1
X_12509_ _05652_ _05605_ VPWR VGND _05664_ sg13g2_nor2b_1
X_12510_ _05663_ _05664_ VPWR VGND _05665_ sg13g2_or2_1
X_12511_ _05665_ VPWR VGND _05666_ sg13g2_buf_1
X_12512_ _05641_ VPWR VGND _05667_ sg13g2_inv_1
X_12513_ _02302_ _05667_ _05656_ _05642_ VPWR VGND 
+ _05668_
+ sg13g2_a22oi_1
X_12514_ _02451_ _05666_ _05668_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[51]\ sg13g2_o21ai_1
X_12515_ _05591_ _05649_ _05660_ VPWR VGND _05669_ sg13g2_a21o_1
X_12516_ _02592_ _05652_ _05669_ _05605_ VPWR VGND 
+ _05670_
+ sg13g2_a22oi_1
X_12517_ _05670_ VPWR VGND _05671_ sg13g2_inv_1
X_12518_ _02302_ _05656_ _05671_ _02450_ VPWR VGND 
+ _05672_
+ sg13g2_a22oi_1
X_12519_ _05657_ _05666_ _05672_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[52]\ sg13g2_o21ai_1
X_12520_ _05642_ _05671_ VPWR VGND _05673_ sg13g2_nand2_1
X_12521_ _02303_ _05666_ _05673_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[53]\ sg13g2_o21ai_1
X_12522_ _03950_ VPWR VGND _05674_ sg13g2_inv_1
X_12523_ _02110_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ _02299_ VPWR VGND 
+ _05675_
+ sg13g2_a22oi_1
X_12524_ _02298_ _02111_ _00081_ VPWR VGND _05676_ sg13g2_or3_1
X_12525_ _00080_ VPWR VGND _05677_ sg13g2_buf_1
X_12526_ _05675_ _05676_ _05677_ VPWR VGND _05678_ sg13g2_a21o_1
X_12527_ _02095_ _05678_ VPWR VGND _05679_ sg13g2_or2_1
X_12528_ _02298_ _02110_ VPWR VGND _05680_ sg13g2_or2_1
X_12529_ _05680_ VPWR VGND _05681_ sg13g2_buf_1
X_12530_ _02111_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _02299_ VPWR VGND 
+ _05682_
+ sg13g2_a22oi_1
X_12531_ _00083_ _05681_ _05682_ VPWR VGND _05683_ sg13g2_o21ai_1
X_12532_ _05683_ VPWR VGND _05684_ sg13g2_buf_1
X_12533_ _02095_ _05684_ _02101_ VPWR VGND _05685_ sg13g2_a21oi_1
X_12534_ _02111_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ _02299_ VPWR VGND 
+ _05686_
+ sg13g2_a22oi_1
X_12535_ _00085_ _05681_ _05686_ VPWR VGND _05687_ sg13g2_o21ai_1
X_12536_ _05687_ VPWR VGND _05688_ sg13g2_buf_1
X_12537_ _02102_ _05688_ VPWR VGND _05689_ sg13g2_nor2_1
X_12538_ _05679_ _05685_ _05689_ _05678_ VPWR VGND 
+ _05690_
+ sg13g2_a22oi_1
X_12539_ _05690_ VPWR VGND _05691_ sg13g2_buf_1
X_12540_ _02299_ _02111_ VPWR VGND _05692_ sg13g2_nor2_1
X_12541_ _02111_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ VPWR VGND _05693_ sg13g2_and2_1
X_12542_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _05692_ _05693_ VPWR VGND _05694_ sg13g2_a21o_1
X_12543_ _02111_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _02299_ VPWR VGND 
+ _05695_
+ sg13g2_a22oi_1
X_12544_ _05695_ VPWR VGND _05696_ sg13g2_buf_1
X_12545_ _02299_ _02111_ _00087_ VPWR VGND _05697_ sg13g2_or3_1
X_12546_ _05697_ VPWR VGND _05698_ sg13g2_buf_1
X_12547_ _02101_ _02094_ VPWR VGND _05699_ sg13g2_or2_1
X_12548_ _05696_ _05698_ _05699_ VPWR VGND _05700_ sg13g2_a21oi_1
X_12549_ _02094_ _05688_ _05694_ _02101_ _05700_ VPWR 
+ VGND
+ _05701_ sg13g2_a221oi_1
X_12550_ _05701_ VPWR VGND _05702_ sg13g2_buf_1
X_12551_ _05702_ VPWR VGND _05703_ sg13g2_inv_1
X_12552_ _02101_ _02094_ VPWR VGND _05704_ sg13g2_nor2_1
X_12553_ _05696_ _05698_ _02102_ VPWR VGND _05705_ sg13g2_a21oi_1
X_12554_ _02094_ _05684_ _05688_ _05704_ _05705_ VPWR 
+ VGND
+ _05706_ sg13g2_a221oi_1
X_12555_ _02105_ _02098_ VPWR VGND _05707_ sg13g2_nor2_1
X_12556_ _05707_ VPWR VGND _05708_ sg13g2_inv_1
X_12557_ _05706_ _05708_ VPWR VGND _05709_ sg13g2_nor2_1
X_12558_ _02098_ _05691_ _05703_ _02105_ _05709_ VPWR 
+ VGND
+ _05710_ sg13g2_a221oi_1
X_12559_ _05710_ VPWR VGND _05711_ sg13g2_buf_1
X_12560_ _05702_ _02098_ VPWR VGND _05712_ sg13g2_nand2b_1
X_12561_ _05696_ _05698_ _02095_ VPWR VGND _05713_ sg13g2_a21oi_1
X_12562_ _05704_ _05694_ _05713_ VPWR VGND _05714_ sg13g2_a21o_1
X_12563_ _05707_ _05714_ VPWR VGND _05715_ sg13g2_nand2_1
X_12564_ _05712_ _05715_ VPWR VGND _05716_ sg13g2_nand2_1
X_12565_ _05702_ _05707_ VPWR VGND _05717_ sg13g2_nand2b_1
X_12566_ _02105_ _05714_ VPWR VGND _05718_ sg13g2_nand2_1
X_12567_ _05706_ _02098_ VPWR VGND _05719_ sg13g2_nand2b_1
X_12568_ _05717_ _05718_ _05719_ VPWR VGND _05720_ sg13g2_nand3_1
X_12569_ _05720_ VPWR VGND _05721_ sg13g2_buf_1
X_12570_ _04119_ _03950_ VPWR VGND _05722_ sg13g2_nor2_1
X_12571_ _04119_ _05716_ _05721_ _05722_ VPWR VGND 
+ _05723_
+ sg13g2_a22oi_1
X_12572_ _05674_ _05711_ _05723_ VPWR VGND _05724_ sg13g2_o21ai_1
X_12573_ _05724_ VPWR VGND _05725_ sg13g2_buf_1
X_12574_ _00082_ VPWR VGND _05726_ sg13g2_inv_1
X_12575_ _05675_ _05676_ VPWR VGND _05727_ sg13g2_and2_1
X_12576_ _05727_ VPWR VGND _05728_ sg13g2_buf_1
X_12577_ _02094_ _05728_ VPWR VGND _05729_ sg13g2_nor2_1
X_12578_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ _02299_ VPWR VGND _05730_ sg13g2_nand2b_1
X_12579_ _02299_ _00079_ VPWR VGND _05731_ sg13g2_nand2b_1
X_12580_ _05730_ _05731_ _02111_ VPWR VGND _05732_ sg13g2_a21oi_1
X_12581_ _02095_ _05677_ _05732_ VPWR VGND _05733_ sg13g2_nor3_1
X_12582_ _02101_ _05729_ _05733_ VPWR VGND _05734_ sg13g2_or3_1
X_12583_ _05734_ VPWR VGND _05735_ sg13g2_buf_1
X_12584_ _02102_ _05684_ VPWR VGND _05736_ sg13g2_nor2_1
X_12585_ _05677_ _05732_ _05736_ VPWR VGND _05737_ sg13g2_o21ai_1
X_12586_ _05737_ VPWR VGND _05738_ sg13g2_buf_1
X_12587_ _02098_ _05726_ _05735_ _05738_ VPWR VGND 
+ _05739_
+ sg13g2_nand4_1
X_12588_ _02099_ _05691_ _02105_ VPWR VGND _05740_ sg13g2_a21oi_1
X_12589_ _02105_ _05706_ VPWR VGND _05741_ sg13g2_and2_1
X_12590_ _05726_ _05735_ _05738_ VPWR VGND _05742_ sg13g2_nand3_1
X_12591_ _05739_ _05740_ _05741_ _05742_ _05674_ VPWR 
+ VGND
+ _05743_ sg13g2_a221oi_1
X_12592_ _04120_ _05721_ VPWR VGND _05744_ sg13g2_nand2_1
X_12593_ _05711_ _05722_ VPWR VGND _05745_ sg13g2_nand2b_1
X_12594_ _05743_ _05744_ _05745_ VPWR VGND _05746_ sg13g2_nand3b_1
X_12595_ _03947_ _03787_ VPWR VGND _05747_ sg13g2_nor2_1
X_12596_ _03947_ _05725_ _05746_ _05747_ VPWR VGND 
+ _05748_
+ sg13g2_a22oi_1
X_12597_ _04120_ _05711_ VPWR VGND _05749_ sg13g2_nand2_1
X_12598_ _04120_ _03950_ VPWR VGND _05750_ sg13g2_nand2b_1
X_12599_ _00084_ VPWR VGND _05751_ sg13g2_buf_1
X_12600_ _05677_ _05732_ _02095_ VPWR VGND _05752_ sg13g2_mux2_1
X_12601_ _02101_ _05677_ VPWR VGND _05753_ sg13g2_and2_1
X_12602_ _05753_ VPWR VGND _05754_ sg13g2_buf_1
X_12603_ _02102_ _05752_ _05754_ _05728_ _00082_ VPWR 
+ VGND
+ _05755_ sg13g2_a221oi_1
X_12604_ _02106_ _05691_ _05755_ VPWR VGND _05756_ sg13g2_nor3_1
X_12605_ _02105_ _02099_ _05755_ VPWR VGND _05757_ sg13g2_nor3_1
X_12606_ _05735_ _05738_ _05708_ VPWR VGND _05758_ sg13g2_a21oi_1
X_12607_ _05751_ _05756_ _05757_ _05758_ VPWR VGND 
+ _05759_
+ sg13g2_nor4_1
X_12608_ _05749_ _05750_ _05759_ VPWR VGND _05760_ sg13g2_a21o_1
X_12609_ _05739_ _05740_ _05741_ _05742_ VPWR VGND 
+ _05761_
+ sg13g2_a22oi_1
X_12610_ _05761_ _05722_ VPWR VGND _05762_ sg13g2_nand2b_1
X_12611_ _03787_ _05760_ _05762_ VPWR VGND _05763_ sg13g2_nand3_1
X_12612_ _05748_ _05763_ VPWR VGND _05764_ sg13g2_and2_1
X_12613_ _05764_ VPWR VGND _05765_ sg13g2_buf_1
X_12614_ _05712_ _05715_ _04119_ VPWR VGND _05766_ sg13g2_a21oi_1
X_12615_ _05721_ _05766_ _05674_ VPWR VGND _05767_ sg13g2_mux2_1
X_12616_ _03787_ _05725_ _05767_ _05747_ VPWR VGND 
+ _05768_
+ sg13g2_a22oi_1
X_12617_ _05768_ VPWR VGND _05769_ sg13g2_inv_1
X_12618_ _03784_ _03605_ VPWR VGND _05770_ sg13g2_nor2_1
X_12619_ _03947_ _05767_ VPWR VGND _05771_ sg13g2_and2_1
X_12620_ _03787_ _05746_ _05747_ _05725_ _05771_ VPWR 
+ VGND
+ _05772_ sg13g2_a221oi_1
X_12621_ _05772_ VPWR VGND _05773_ sg13g2_inv_1
X_12622_ _03784_ _05769_ _05770_ _05773_ VPWR VGND 
+ _05774_
+ sg13g2_a22oi_1
X_12623_ _03606_ _05765_ _05774_ VPWR VGND _05775_ sg13g2_o21ai_1
X_12624_ _02771_ _05770_ VPWR VGND _05776_ sg13g2_nand2_1
X_12625_ _05696_ _05698_ VPWR VGND _05777_ sg13g2_nand2_1
X_12626_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ _05547_ _05777_ VPWR VGND _05778_ sg13g2_nor3_1
X_12627_ _05564_ _05702_ _05778_ VPWR VGND _05779_ sg13g2_nand3_1
X_12628_ _05570_ _05721_ _05725_ _05779_ VPWR VGND 
+ _05780_
+ sg13g2_nor4_1
X_12629_ _05768_ _05776_ _05780_ VPWR VGND _05781_ sg13g2_o21ai_1
X_12630_ _05781_ _05632_ _05772_ VPWR VGND _05782_ sg13g2_nand3b_1
X_12631_ _05775_ _05782_ VPWR VGND _05783_ sg13g2_nor2_1
X_12632_ _05744_ _05745_ VPWR VGND _05784_ sg13g2_nand2_1
X_12633_ _05743_ _05784_ VPWR VGND _05785_ sg13g2_nor2_1
X_12634_ _00086_ VPWR VGND _05786_ sg13g2_inv_1
X_12635_ _02099_ _00082_ VPWR VGND _05787_ sg13g2_nor2_1
X_12636_ _02102_ _05752_ _05754_ _05728_ _02098_ VPWR 
+ VGND
+ _05788_ sg13g2_a221oi_1
X_12637_ _02105_ _05787_ _05788_ VPWR VGND _05789_ sg13g2_or3_1
X_12638_ _05789_ VPWR VGND _05790_ sg13g2_buf_1
X_12639_ _02105_ _00082_ VPWR VGND _05791_ sg13g2_nand2_1
X_12640_ _05735_ _05738_ _05791_ VPWR VGND _05792_ sg13g2_a21o_1
X_12641_ _05751_ _05790_ _05792_ VPWR VGND _05793_ sg13g2_nand3b_1
X_12642_ _05761_ _05793_ _04120_ VPWR VGND _05794_ sg13g2_nand3b_1
X_12643_ _05756_ _05757_ _05758_ VPWR VGND _05795_ sg13g2_or3_1
X_12644_ _05795_ VPWR VGND _05796_ sg13g2_buf_1
X_12645_ _04120_ _05674_ VPWR VGND _05797_ sg13g2_nor2_1
X_12646_ _05722_ _05796_ _05797_ _05793_ VPWR VGND 
+ _05798_
+ sg13g2_a22oi_1
X_12647_ _05786_ _05794_ _05798_ VPWR VGND _05799_ sg13g2_nand3_1
X_12648_ _03947_ _05785_ _05799_ VPWR VGND _05800_ sg13g2_nand3_1
X_12649_ _03947_ VPWR VGND _05801_ sg13g2_inv_1
X_12650_ _05801_ _03787_ VPWR VGND _05802_ sg13g2_nand2_1
X_12651_ _05802_ _05799_ VPWR VGND _05803_ sg13g2_nand2b_1
X_12652_ _05760_ _05762_ VPWR VGND _05804_ sg13g2_nand2_1
X_12653_ _05747_ _05804_ VPWR VGND _05805_ sg13g2_nand2_1
X_12654_ _05800_ _05803_ _05805_ VPWR VGND _05806_ sg13g2_nand3_1
X_12655_ _05765_ VPWR VGND _05807_ sg13g2_inv_1
X_12656_ _03784_ _05773_ _05770_ _05807_ VPWR VGND 
+ _05808_
+ sg13g2_a22oi_1
X_12657_ _03606_ _05806_ _05808_ VPWR VGND _05809_ sg13g2_o21ai_1
X_12658_ _01901_ _05809_ _05652_ VPWR VGND _05810_ sg13g2_a21oi_1
X_12659_ _05666_ _05783_ _05810_ VPWR VGND _05811_ sg13g2_and3_1
X_12660_ _00088_ VPWR VGND _05812_ sg13g2_inv_1
X_12661_ _05794_ _05798_ VPWR VGND _05813_ sg13g2_nand2_1
X_12662_ _05747_ _05813_ VPWR VGND _05814_ sg13g2_and2_1
X_12663_ _05674_ _05790_ _05792_ VPWR VGND _05815_ sg13g2_nand3_1
X_12664_ _05674_ _05751_ _05815_ VPWR VGND _05816_ sg13g2_o21ai_1
X_12665_ _05751_ _05796_ VPWR VGND _05817_ sg13g2_nand2_1
X_12666_ _05816_ _05817_ _04120_ VPWR VGND _05818_ sg13g2_mux2_1
X_12667_ _05760_ _05762_ _05801_ VPWR VGND _05819_ sg13g2_a21o_1
X_12668_ _05786_ _05818_ _05819_ _05802_ VPWR VGND 
+ _05820_
+ sg13g2_a22oi_1
X_12669_ _05814_ _05820_ VPWR VGND _05821_ sg13g2_nor2_1
X_12670_ _03784_ _05765_ VPWR VGND _05822_ sg13g2_nand2_1
X_12671_ _03785_ _03605_ VPWR VGND _05823_ sg13g2_nand2_1
X_12672_ _05812_ _05821_ _05822_ _05823_ VPWR VGND 
+ _05824_
+ sg13g2_a22oi_1
X_12673_ _05770_ _05806_ _05824_ VPWR VGND _05825_ sg13g2_a21oi_1
X_12674_ _01901_ _05825_ VPWR VGND _05826_ sg13g2_nand2_1
X_12675_ _02759_ _05623_ _02766_ VPWR VGND _05827_ sg13g2_a21o_1
X_12676_ _05575_ _05578_ VPWR VGND _05828_ sg13g2_nor2_1
X_12677_ _02094_ _05684_ _05705_ VPWR VGND _05829_ sg13g2_a21oi_1
X_12678_ _03591_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _05531_ _05688_ VPWR VGND 
+ _05830_
+ sg13g2_nor4_1
X_12679_ _05550_ _05829_ _05711_ _05830_ VPWR VGND 
+ _05831_
+ sg13g2_nand4_1
X_12680_ _02926_ _05572_ VPWR VGND _05832_ sg13g2_nor2_1
X_12681_ _05571_ _05832_ _05765_ VPWR VGND _05833_ sg13g2_o21ai_1
X_12682_ _05828_ _05746_ _05831_ _05833_ VPWR VGND 
+ _05834_
+ sg13g2_or4_1
X_12683_ _02771_ _05775_ _05827_ _05633_ _05834_ VPWR 
+ VGND
+ _05835_ sg13g2_a221oi_1
X_12684_ _05809_ _05835_ VPWR VGND _05836_ sg13g2_nor2b_1
X_12685_ _05656_ _05826_ _05836_ VPWR VGND _05837_ sg13g2_nand3b_1
X_12686_ _03787_ _05725_ VPWR VGND _05838_ sg13g2_and2_1
X_12687_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _05568_ _05693_ _05714_ VPWR VGND 
+ _05839_
+ sg13g2_nor4_1
X_12688_ _05712_ _05839_ VPWR VGND _05840_ sg13g2_nand2_1
X_12689_ _05626_ _05838_ _05767_ _05840_ VPWR VGND 
+ _05841_
+ sg13g2_nor4_1
X_12690_ _03605_ _05773_ _05649_ VPWR VGND _05842_ sg13g2_a21oi_1
X_12691_ _01901_ _05775_ _05669_ VPWR VGND _05843_ sg13g2_a21oi_1
X_12692_ _05670_ _05841_ _05842_ _05843_ VPWR VGND 
+ _05844_
+ sg13g2_and4_1
X_12693_ _05844_ VPWR VGND _05845_ sg13g2_inv_1
X_12694_ _05811_ _05837_ _05845_ VPWR VGND _05846_ sg13g2_a21oi_1
X_12695_ _04120_ _05751_ _05796_ VPWR VGND _05847_ sg13g2_nand3_1
X_12696_ _04120_ _05816_ _05847_ VPWR VGND _05848_ sg13g2_o21ai_1
X_12697_ _05848_ _00086_ _03787_ VPWR VGND _05849_ sg13g2_mux2_1
X_12698_ _05801_ _05786_ VPWR VGND _05850_ sg13g2_nor2_1
X_12699_ _05801_ _05849_ _05850_ _05813_ _03605_ VPWR 
+ VGND
+ _05851_ sg13g2_a221oi_1
X_12700_ _03605_ _05812_ _05851_ VPWR VGND _05852_ sg13g2_a21oi_1
X_12701_ _03785_ _05812_ VPWR VGND _05853_ sg13g2_nor2_1
X_12702_ _05814_ _05820_ VPWR VGND _05854_ sg13g2_or2_1
X_12703_ _03785_ _05852_ _05853_ _05854_ VPWR VGND 
+ _05855_
+ sg13g2_a22oi_1
X_12704_ _00089_ VPWR VGND _05856_ sg13g2_inv_1
X_12705_ _02771_ _01901_ VPWR VGND _05857_ sg13g2_nor2_1
X_12706_ _02771_ _05825_ _05855_ _05856_ _05857_ VPWR 
+ VGND
+ _05858_ sg13g2_a221oi_1
X_12707_ _05800_ _05803_ _05805_ VPWR VGND _05859_ sg13g2_and3_1
X_12708_ _05801_ _05849_ _05850_ _05813_ _00088_ VPWR 
+ VGND
+ _05860_ sg13g2_a221oi_1
X_12709_ _05859_ _05860_ VPWR VGND _05861_ sg13g2_nor2_1
X_12710_ _05823_ _05860_ VPWR VGND _05862_ sg13g2_nor2_1
X_12711_ _05770_ _05854_ _05861_ _03784_ _05862_ VPWR 
+ VGND
+ _05863_ sg13g2_a221oi_1
X_12712_ _05500_ _05501_ _05675_ _05681_ _00081_ VPWR 
+ VGND
+ _05864_ sg13g2_a221oi_1
X_12713_ _05498_ _05561_ VPWR VGND _05865_ sg13g2_nor2_1
X_12714_ _05496_ _05508_ _05865_ VPWR VGND _05866_ sg13g2_o21ai_1
X_12715_ _05735_ _05738_ _05864_ _05866_ VPWR VGND 
+ _05867_
+ sg13g2_nand4_1
X_12716_ _05584_ _05796_ _05867_ VPWR VGND _05868_ sg13g2_or3_1
X_12717_ _05609_ _05813_ _05820_ _05868_ VPWR VGND 
+ _05869_
+ sg13g2_nor4_1
X_12718_ _05607_ _05614_ _05863_ _05869_ VPWR VGND 
+ _05870_
+ sg13g2_nand4_1
X_12719_ _05858_ _05870_ VPWR VGND _05871_ sg13g2_nor2_1
X_12720_ _03264_ _05504_ VPWR VGND _05872_ sg13g2_nand2_1
X_12721_ _03415_ _05872_ VPWR VGND _05873_ sg13g2_nor2_1
X_12722_ _03415_ _05504_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2931_o\ VPWR VGND _05874_ sg13g2_a21oi_1
X_12723_ _03591_ _05874_ _05684_ VPWR VGND _05875_ sg13g2_o21ai_1
X_12724_ _00083_ _05873_ _05875_ VPWR VGND _05876_ sg13g2_nor3_1
X_12725_ _05576_ _05691_ _05876_ VPWR VGND _05877_ sg13g2_and3_1
X_12726_ _05583_ _05586_ VPWR VGND _05878_ sg13g2_nor2_1
X_12727_ _05878_ _05804_ VPWR VGND _05879_ sg13g2_nor2_1
X_12728_ _05558_ _05761_ _05877_ _05879_ VPWR VGND 
+ _05880_
+ sg13g2_nand4_1
X_12729_ _05595_ _05806_ _05824_ _05880_ VPWR VGND 
+ _05881_
+ sg13g2_or4_1
X_12730_ _02771_ _05809_ _05863_ _05856_ _05857_ VPWR 
+ VGND
+ _05882_ sg13g2_a221oi_1
X_12731_ _05641_ _05881_ _05882_ VPWR VGND _05883_ sg13g2_or3_1
X_12732_ _05786_ _05747_ VPWR VGND _05884_ sg13g2_nor2_1
X_12733_ _05801_ _05813_ _05884_ VPWR VGND _05885_ sg13g2_o21ai_1
X_12734_ _05790_ _05792_ VPWR VGND _05886_ sg13g2_nand2_1
X_12735_ _02102_ _05752_ _05754_ _05728_ VPWR VGND 
+ _05887_
+ sg13g2_a22oi_1
X_12736_ _00079_ _05514_ _05732_ VPWR VGND _05888_ sg13g2_nor3_1
X_12737_ _05517_ _05887_ _05888_ VPWR VGND _05889_ sg13g2_nand3b_1
X_12738_ _05556_ _05584_ VPWR VGND _05890_ sg13g2_nor2_1
X_12739_ _05557_ _05587_ _05890_ VPWR VGND _05891_ sg13g2_nor3_1
X_12740_ _05886_ _05848_ _05889_ _05891_ VPWR VGND 
+ _05892_
+ sg13g2_nor4_1
X_12741_ _05604_ _05885_ _05892_ VPWR VGND _05893_ sg13g2_nand3_1
X_12742_ _02596_ _02592_ _00076_ VPWR VGND _05894_ sg13g2_o21ai_1
X_12743_ _02596_ _05614_ _05894_ VPWR VGND _05895_ sg13g2_a21oi_1
X_12744_ _05893_ _05895_ VPWR VGND _05896_ sg13g2_nor2_1
X_12745_ _02771_ _01901_ _00089_ VPWR VGND _05897_ sg13g2_o21ai_1
X_12746_ _02771_ _05863_ _05897_ VPWR VGND _05898_ sg13g2_a21o_1
X_12747_ _05855_ _05896_ _05898_ VPWR VGND _05899_ sg13g2_nand3_1
X_12748_ _05871_ _05883_ _05899_ VPWR VGND _05900_ sg13g2_a21oi_1
X_12749_ _05846_ _05900_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[0]\ sg13g2_xor2_1
X_12750_ _05846_ _05900_ VPWR VGND _05901_ sg13g2_or2_1
X_12751_ _05899_ _05871_ VPWR VGND _05902_ sg13g2_nand2b_1
X_12752_ _05844_ _05811_ VPWR VGND _05903_ sg13g2_nand2_1
X_12753_ _05902_ _05903_ VPWR VGND _05904_ sg13g2_xor2_1
X_12754_ _05901_ _05904_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[1]\ sg13g2_xnor2_1
X_12755_ _05902_ _05903_ VPWR VGND _05905_ sg13g2_nand2_1
X_12756_ _05902_ _05903_ VPWR VGND _05906_ sg13g2_nor2_1
X_12757_ _05901_ _05905_ _05906_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[2]\ sg13g2_a21oi_1
X_12758_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2463_q\ _01102_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1321_o\ sg13g2_nand2b_1
X_12759_ _05469_ _04331_ VPWR VGND _05907_ sg13g2_nor2_1
X_12760_ _05469_ _05069_ _05907_ VPWR VGND \atbs_core_0.dac_control_0.n1498_o\ sg13g2_a21oi_1
X_12761_ \atbs_core_0.dac_control_0.n1592_q[0]\ \atbs_core_0.dac_control_0.dac_counter_strb\ VPWR VGND \atbs_core_0.dac_control_0.n1566_o[0]\ sg13g2_nor2_1
X_12762_ \atbs_core_0.dac_control_0.n1592_q[1]\ \atbs_core_0.dac_control_0.n1592_q[0]\ VPWR VGND _05908_ sg13g2_xnor2_1
X_12763_ \atbs_core_0.dac_control_0.dac_counter_strb\ _05908_ VPWR VGND \atbs_core_0.dac_control_0.n1566_o[1]\ sg13g2_nor2_1
X_12764_ _00030_ _04620_ VPWR VGND _05909_ sg13g2_xnor2_1
X_12765_ \atbs_core_0.dac_control_0.dac_counter_strb\ _05909_ VPWR VGND \atbs_core_0.dac_control_0.n1566_o[2]\ sg13g2_nor2_1
X_12766_ \atbs_core_0.dac_control_1.n1727_q[0]\ \atbs_core_0.dac_control_1.dac_counter_strb\ VPWR VGND \atbs_core_0.dac_control_1.n1701_o[0]\ sg13g2_nor2_1
X_12767_ \atbs_core_0.dac_control_1.n1727_q[1]\ \atbs_core_0.dac_control_1.n1727_q[0]\ VPWR VGND _05910_ sg13g2_xnor2_1
X_12768_ \atbs_core_0.dac_control_1.dac_counter_strb\ _05910_ VPWR VGND \atbs_core_0.dac_control_1.n1701_o[1]\ sg13g2_nor2_1
X_12769_ _00053_ _04828_ VPWR VGND _05911_ sg13g2_xnor2_1
X_12770_ \atbs_core_0.dac_control_1.dac_counter_strb\ _05911_ VPWR VGND \atbs_core_0.dac_control_1.n1701_o[2]\ sg13g2_nor2_1
X_12771_ _04831_ _04830_ VPWR VGND _05912_ sg13g2_or2_1
X_12772_ \atbs_core_0.debouncer_0.bouncing_sync\ _04837_ VPWR VGND _05913_ sg13g2_xnor2_1
X_12773_ _05912_ _05913_ _04836_ VPWR VGND _05914_ sg13g2_o21ai_1
X_12774_ _05914_ VPWR VGND _05915_ sg13g2_buf_1
X_12775_ _04833_ _05915_ VPWR VGND \atbs_core_0.debouncer_0.n1128_o[0]\ sg13g2_nor2_1
X_12776_ _04833_ _04832_ VPWR VGND _05916_ sg13g2_xnor2_1
X_12777_ _05915_ _05916_ VPWR VGND \atbs_core_0.debouncer_0.n1128_o[1]\ sg13g2_nor2_1
X_12778_ _04833_ _04832_ VPWR VGND _05917_ sg13g2_nand2_1
X_12779_ \atbs_core_0.debouncer_0.counter_value[2]\ _05917_ VPWR VGND _05918_ sg13g2_xor2_1
X_12780_ _05915_ _05918_ VPWR VGND \atbs_core_0.debouncer_0.n1128_o[2]\ sg13g2_nor2_1
X_12781_ _04833_ _04832_ \atbs_core_0.debouncer_0.counter_value[2]\ VPWR VGND _05919_ sg13g2_nand3_1
X_12782_ \atbs_core_0.debouncer_0.counter_value[3]\ _05919_ VPWR VGND _05920_ sg13g2_xor2_1
X_12783_ _05915_ _05920_ VPWR VGND \atbs_core_0.debouncer_0.n1128_o[3]\ sg13g2_nor2_1
X_12784_ _04847_ _04846_ VPWR VGND _05921_ sg13g2_or2_1
X_12785_ \atbs_core_0.debouncer_1.bouncing_sync\ _04853_ VPWR VGND _05922_ sg13g2_xnor2_1
X_12786_ _05921_ _05922_ _04852_ VPWR VGND _05923_ sg13g2_o21ai_1
X_12787_ _05923_ VPWR VGND _05924_ sg13g2_buf_1
X_12788_ _04849_ _05924_ VPWR VGND \atbs_core_0.debouncer_1.n1128_o[0]\ sg13g2_nor2_1
X_12789_ _04849_ _04848_ VPWR VGND _05925_ sg13g2_xnor2_1
X_12790_ _05924_ _05925_ VPWR VGND \atbs_core_0.debouncer_1.n1128_o[1]\ sg13g2_nor2_1
X_12791_ _04849_ _04848_ VPWR VGND _05926_ sg13g2_nand2_1
X_12792_ \atbs_core_0.debouncer_1.counter_value[2]\ _05926_ VPWR VGND _05927_ sg13g2_xor2_1
X_12793_ _05924_ _05927_ VPWR VGND \atbs_core_0.debouncer_1.n1128_o[2]\ sg13g2_nor2_1
X_12794_ _04849_ _04848_ \atbs_core_0.debouncer_1.counter_value[2]\ VPWR VGND _05928_ sg13g2_nand3_1
X_12795_ \atbs_core_0.debouncer_1.counter_value[3]\ _05928_ VPWR VGND _05929_ sg13g2_xor2_1
X_12796_ _05924_ _05929_ VPWR VGND \atbs_core_0.debouncer_1.n1128_o[3]\ sg13g2_nor2_1
X_12797_ _04863_ _04862_ VPWR VGND _05930_ sg13g2_or2_1
X_12798_ \atbs_core_0.debouncer_2.bouncing_sync\ _04869_ VPWR VGND _05931_ sg13g2_xnor2_1
X_12799_ _05930_ _05931_ _04868_ VPWR VGND _05932_ sg13g2_o21ai_1
X_12800_ _05932_ VPWR VGND _05933_ sg13g2_buf_1
X_12801_ _04865_ _05933_ VPWR VGND \atbs_core_0.debouncer_2.n1128_o[0]\ sg13g2_nor2_1
X_12802_ _04865_ _04864_ VPWR VGND _05934_ sg13g2_xnor2_1
X_12803_ _05933_ _05934_ VPWR VGND \atbs_core_0.debouncer_2.n1128_o[1]\ sg13g2_nor2_1
X_12804_ _04865_ _04864_ VPWR VGND _05935_ sg13g2_nand2_1
X_12805_ \atbs_core_0.debouncer_2.counter_value[2]\ _05935_ VPWR VGND _05936_ sg13g2_xor2_1
X_12806_ _05933_ _05936_ VPWR VGND \atbs_core_0.debouncer_2.n1128_o[2]\ sg13g2_nor2_1
X_12807_ _04865_ _04864_ \atbs_core_0.debouncer_2.counter_value[2]\ VPWR VGND _05937_ sg13g2_nand3_1
X_12808_ \atbs_core_0.debouncer_2.counter_value[3]\ _05937_ VPWR VGND _05938_ sg13g2_xor2_1
X_12809_ _05933_ _05938_ VPWR VGND \atbs_core_0.debouncer_2.n1128_o[3]\ sg13g2_nor2_1
X_12810_ _04878_ _04879_ VPWR VGND _05939_ sg13g2_or2_1
X_12811_ \atbs_core_0.debouncer_3.bouncing_sync\ _04885_ VPWR VGND _05940_ sg13g2_xnor2_1
X_12812_ _05939_ _05940_ _04884_ VPWR VGND _05941_ sg13g2_o21ai_1
X_12813_ _05941_ VPWR VGND _05942_ sg13g2_buf_1
X_12814_ _04881_ _05942_ VPWR VGND \atbs_core_0.debouncer_3.n1128_o[0]\ sg13g2_nor2_1
X_12815_ _04881_ _04880_ VPWR VGND _05943_ sg13g2_xnor2_1
X_12816_ _05942_ _05943_ VPWR VGND \atbs_core_0.debouncer_3.n1128_o[1]\ sg13g2_nor2_1
X_12817_ _04881_ _04880_ VPWR VGND _05944_ sg13g2_nand2_1
X_12818_ \atbs_core_0.debouncer_3.counter_value[2]\ _05944_ VPWR VGND _05945_ sg13g2_xor2_1
X_12819_ _05942_ _05945_ VPWR VGND \atbs_core_0.debouncer_3.n1128_o[2]\ sg13g2_nor2_1
X_12820_ _04881_ _04880_ \atbs_core_0.debouncer_3.counter_value[2]\ VPWR VGND _05946_ sg13g2_nand3_1
X_12821_ \atbs_core_0.debouncer_3.counter_value[3]\ _05946_ VPWR VGND _05947_ sg13g2_xor2_1
X_12822_ _05942_ _05947_ VPWR VGND \atbs_core_0.debouncer_3.n1128_o[3]\ sg13g2_nor2_1
X_12823_ _04895_ _04894_ VPWR VGND _05948_ sg13g2_or2_1
X_12824_ \atbs_core_0.debouncer_4.bouncing_sync\ _04901_ VPWR VGND _05949_ sg13g2_xnor2_1
X_12825_ _05948_ _05949_ _04900_ VPWR VGND _05950_ sg13g2_o21ai_1
X_12826_ _05950_ VPWR VGND _05951_ sg13g2_buf_1
X_12827_ _04897_ _05951_ VPWR VGND \atbs_core_0.debouncer_4.n1128_o[0]\ sg13g2_nor2_1
X_12828_ _04897_ _04896_ VPWR VGND _05952_ sg13g2_xnor2_1
X_12829_ _05951_ _05952_ VPWR VGND \atbs_core_0.debouncer_4.n1128_o[1]\ sg13g2_nor2_1
X_12830_ _04897_ _04896_ VPWR VGND _05953_ sg13g2_nand2_1
X_12831_ \atbs_core_0.debouncer_4.counter_value[2]\ _05953_ VPWR VGND _05954_ sg13g2_xor2_1
X_12832_ _05951_ _05954_ VPWR VGND \atbs_core_0.debouncer_4.n1128_o[2]\ sg13g2_nor2_1
X_12833_ _04897_ _04896_ \atbs_core_0.debouncer_4.counter_value[2]\ VPWR VGND _05955_ sg13g2_nand3_1
X_12834_ \atbs_core_0.debouncer_4.counter_value[3]\ _05955_ VPWR VGND _05956_ sg13g2_xor2_1
X_12835_ _05951_ _05956_ VPWR VGND \atbs_core_0.debouncer_4.n1128_o[3]\ sg13g2_nor2_1
X_12836_ _04911_ _04910_ VPWR VGND _05957_ sg13g2_or2_1
X_12837_ \atbs_core_0.debouncer_5.bouncing_sync\ _04917_ VPWR VGND _05958_ sg13g2_xnor2_1
X_12838_ _05957_ _05958_ _04916_ VPWR VGND _05959_ sg13g2_o21ai_1
X_12839_ _05959_ VPWR VGND _05960_ sg13g2_buf_1
X_12840_ _04913_ _05960_ VPWR VGND \atbs_core_0.debouncer_5.n1128_o[0]\ sg13g2_nor2_1
X_12841_ _04913_ _04912_ VPWR VGND _05961_ sg13g2_xnor2_1
X_12842_ _05960_ _05961_ VPWR VGND \atbs_core_0.debouncer_5.n1128_o[1]\ sg13g2_nor2_1
X_12843_ _04913_ _04912_ VPWR VGND _05962_ sg13g2_nand2_1
X_12844_ \atbs_core_0.debouncer_5.counter_value[2]\ _05962_ VPWR VGND _05963_ sg13g2_xor2_1
X_12845_ _05960_ _05963_ VPWR VGND \atbs_core_0.debouncer_5.n1128_o[2]\ sg13g2_nor2_1
X_12846_ _04913_ _04912_ \atbs_core_0.debouncer_5.counter_value[2]\ VPWR VGND _05964_ sg13g2_nand3_1
X_12847_ \atbs_core_0.debouncer_5.counter_value[3]\ _05964_ VPWR VGND _05965_ sg13g2_xor2_1
X_12848_ _05960_ _05965_ VPWR VGND \atbs_core_0.debouncer_5.n1128_o[3]\ sg13g2_nor2_1
X_12849_ _04355_ dac_upper_o[2] dac_upper_o[1] \atbs_core_0.n1068_q[1]\ VPWR VGND 
+ _05966_
+ sg13g2_a22oi_1
X_12850_ _04355_ dac_upper_o[2] \atbs_core_0.n1068_q[3]\ VPWR VGND _05967_ sg13g2_o21ai_1
X_12851_ _04355_ dac_upper_o[3] VPWR VGND _05968_ sg13g2_nand2_1
X_12852_ dac_upper_o[1] dac_upper_o[0] _04343_ VPWR VGND _05969_ sg13g2_a21oi_1
X_12853_ _04343_ _05966_ _05967_ _05968_ _05969_ VPWR 
+ VGND
+ _05970_ sg13g2_a221oi_1
X_12854_ \atbs_core_0.n1068_q[3]\ dac_upper_o[3] _05970_ VPWR VGND _05971_ sg13g2_a21o_1
X_12855_ dac_upper_o[3] dac_upper_o[2] VPWR VGND _05972_ sg13g2_and2_1
X_12856_ _04343_ _05966_ _05969_ VPWR VGND _05973_ sg13g2_a21oi_1
X_12857_ _04343_ _05971_ _05972_ _05973_ VPWR VGND 
+ _05974_
+ sg13g2_a22oi_1
X_12858_ _00078_ _05974_ VPWR VGND _05975_ sg13g2_nand2_1
X_12859_ \atbs_core_0.n1068_q[4]\ dac_upper_o[5] _05975_ VPWR VGND _05976_ sg13g2_and3_1
X_12860_ \atbs_core_0.n1068_q[5]\ _05976_ _04343_ VPWR VGND _05977_ sg13g2_o21ai_1
X_12861_ _00078_ _05974_ VPWR VGND _05978_ sg13g2_nor2_1
X_12862_ \atbs_core_0.n1068_q[4]\ _05978_ _05975_ VPWR VGND _05979_ sg13g2_o21ai_1
X_12863_ dac_upper_o[5] _05979_ VPWR VGND _05980_ sg13g2_nor2b_1
X_12864_ dac_upper_o[1] dac_upper_o[0] dac_upper_o[4] _05972_ VPWR VGND 
+ _05981_
+ sg13g2_and4_1
X_12865_ _05978_ _05981_ dac_upper_o[5] VPWR VGND _05982_ sg13g2_o21ai_1
X_12866_ _05977_ _05980_ _05982_ VPWR VGND _05983_ sg13g2_o21ai_1
X_12867_ dac_upper_o[6] dac_upper_o[7] _05983_ VPWR VGND \atbs_core_0.n148_o\ sg13g2_nand3_1
X_12868_ dac_lower_o[5] dac_lower_o[4] dac_lower_o[7] dac_lower_o[6] VPWR VGND 
+ _05984_
+ sg13g2_nor4_1
X_12869_ dac_lower_o[1] dac_lower_o[0] dac_lower_o[3] dac_lower_o[2] VPWR VGND 
+ _05985_
+ sg13g2_nor4_1
X_12870_ _05984_ _05985_ VPWR VGND \atbs_core_0.n156_o\ sg13g2_nand2_1
X_12871_ _01035_ _01068_ VPWR VGND _05986_ sg13g2_and2_1
X_12872_ _05986_ VPWR VGND _05987_ sg13g2_buf_1
X_12873_ _01071_ _00842_ _01183_ _05987_ VPWR VGND 
+ _05988_
+ sg13g2_nand4_1
X_12874_ \atbs_core_0.main_counter_value[7]\ VPWR VGND _05989_ sg13g2_inv_1
X_12875_ _00835_ _00846_ \atbs_core_0.main_counter_value[2]\ VPWR VGND _05990_ sg13g2_nand3_1
X_12876_ _00847_ _05990_ VPWR VGND _05991_ sg13g2_nor2_1
X_12877_ _00848_ _05991_ VPWR VGND _05992_ sg13g2_and2_1
X_12878_ _05992_ VPWR VGND _05993_ sg13g2_buf_1
X_12879_ _00825_ \atbs_core_0.main_counter_value[6]\ _05993_ VPWR VGND _05994_ sg13g2_nand3_1
X_12880_ _05989_ _05994_ VPWR VGND _05995_ sg13g2_nor2_1
X_12881_ _00836_ _00837_ _00838_ _00833_ VPWR VGND 
+ _05996_
+ sg13g2_and4_1
X_12882_ \atbs_core_0.main_counter_value[19]\ _00832_ _05995_ _05996_ VPWR VGND 
+ _05997_
+ sg13g2_nand4_1
X_12883_ _05071_ _05481_ _05988_ _05997_ VPWR VGND 
+ _05998_
+ sg13g2_nand4_1
X_12884_ _05998_ VPWR VGND _05999_ sg13g2_buf_1
X_12885_ _05999_ VPWR VGND _06000_ sg13g2_buf_1
X_12886_ _00835_ _06000_ VPWR VGND \atbs_core_0.n206_o[0]\ sg13g2_nor2_1
X_12887_ _00827_ _00828_ _05995_ VPWR VGND _06001_ sg13g2_nand3_1
X_12888_ _00836_ _06001_ VPWR VGND _06002_ sg13g2_xor2_1
X_12889_ _06000_ _06002_ VPWR VGND \atbs_core_0.n206_o[10]\ sg13g2_nor2_1
X_12890_ \atbs_core_0.main_counter_value[11]\ VPWR VGND _06003_ sg13g2_inv_1
X_12891_ _00827_ _00828_ _00836_ _05995_ VPWR VGND 
+ _06004_
+ sg13g2_nand4_1
X_12892_ _06003_ _06004_ VPWR VGND _06005_ sg13g2_xnor2_1
X_12893_ _06000_ _06005_ VPWR VGND \atbs_core_0.n206_o[11]\ sg13g2_nor2_1
X_12894_ _06003_ _06004_ VPWR VGND _06006_ sg13g2_nor2_1
X_12895_ _00838_ _06006_ VPWR VGND _06007_ sg13g2_xnor2_1
X_12896_ _06000_ _06007_ VPWR VGND \atbs_core_0.n206_o[12]\ sg13g2_nor2_1
X_12897_ _00838_ _06006_ VPWR VGND _06008_ sg13g2_nand2_1
X_12898_ _00837_ _06008_ VPWR VGND _06009_ sg13g2_xor2_1
X_12899_ _06000_ _06009_ VPWR VGND \atbs_core_0.n206_o[13]\ sg13g2_nor2_1
X_12900_ _00837_ _00838_ _06006_ VPWR VGND _06010_ sg13g2_nand3_1
X_12901_ \atbs_core_0.main_counter_value[14]\ _06010_ VPWR VGND _06011_ sg13g2_xor2_1
X_12902_ _06000_ _06011_ VPWR VGND \atbs_core_0.n206_o[14]\ sg13g2_nor2_1
X_12903_ \atbs_core_0.main_counter_value[15]\ VPWR VGND _06012_ sg13g2_inv_1
X_12904_ _00837_ _00838_ \atbs_core_0.main_counter_value[14]\ _06006_ VPWR VGND 
+ _06013_
+ sg13g2_nand4_1
X_12905_ _06012_ _06013_ VPWR VGND _06014_ sg13g2_xnor2_1
X_12906_ _06000_ _06014_ VPWR VGND \atbs_core_0.n206_o[15]\ sg13g2_nor2_1
X_12907_ _06012_ _06013_ VPWR VGND _06015_ sg13g2_nor2_1
X_12908_ _00830_ _06015_ VPWR VGND _06016_ sg13g2_xnor2_1
X_12909_ _06000_ _06016_ VPWR VGND \atbs_core_0.n206_o[16]\ sg13g2_nor2_1
X_12910_ _00830_ _06015_ VPWR VGND _06017_ sg13g2_nand2_1
X_12911_ _00829_ _06017_ VPWR VGND _06018_ sg13g2_xor2_1
X_12912_ _06000_ _06018_ VPWR VGND \atbs_core_0.n206_o[17]\ sg13g2_nor2_1
X_12913_ _00829_ _00830_ _06015_ VPWR VGND _06019_ sg13g2_nand3_1
X_12914_ _00833_ _06019_ VPWR VGND _06020_ sg13g2_xor2_1
X_12915_ _06000_ _06020_ VPWR VGND \atbs_core_0.n206_o[18]\ sg13g2_nor2_1
X_12916_ _05999_ VPWR VGND _06021_ sg13g2_buf_1
X_12917_ _00829_ _00830_ _00833_ _06015_ VPWR VGND 
+ _06022_
+ sg13g2_nand4_1
X_12918_ \atbs_core_0.main_counter_value[19]\ _06022_ VPWR VGND _06023_ sg13g2_xor2_1
X_12919_ _06021_ _06023_ VPWR VGND \atbs_core_0.n206_o[19]\ sg13g2_nor2_1
X_12920_ _00835_ _00846_ VPWR VGND _06024_ sg13g2_xnor2_1
X_12921_ _06021_ _06024_ VPWR VGND \atbs_core_0.n206_o[1]\ sg13g2_nor2_1
X_12922_ _00835_ _00846_ VPWR VGND _06025_ sg13g2_nand2_1
X_12923_ \atbs_core_0.main_counter_value[2]\ _06025_ VPWR VGND _06026_ sg13g2_xor2_1
X_12924_ _06021_ _06026_ VPWR VGND \atbs_core_0.n206_o[2]\ sg13g2_nor2_1
X_12925_ _00847_ _05990_ VPWR VGND _06027_ sg13g2_xnor2_1
X_12926_ _06021_ _06027_ VPWR VGND \atbs_core_0.n206_o[3]\ sg13g2_nor2_1
X_12927_ _00848_ _05991_ VPWR VGND _06028_ sg13g2_xnor2_1
X_12928_ _06021_ _06028_ VPWR VGND \atbs_core_0.n206_o[4]\ sg13g2_nor2_1
X_12929_ _00825_ _05993_ VPWR VGND _06029_ sg13g2_xnor2_1
X_12930_ _06021_ _06029_ VPWR VGND \atbs_core_0.n206_o[5]\ sg13g2_nor2_1
X_12931_ _00825_ _05993_ VPWR VGND _06030_ sg13g2_nand2_1
X_12932_ \atbs_core_0.main_counter_value[6]\ _06030_ VPWR VGND _06031_ sg13g2_xor2_1
X_12933_ _06021_ _06031_ VPWR VGND \atbs_core_0.n206_o[6]\ sg13g2_nor2_1
X_12934_ _05989_ _05994_ VPWR VGND _06032_ sg13g2_xnor2_1
X_12935_ _06021_ _06032_ VPWR VGND \atbs_core_0.n206_o[7]\ sg13g2_nor2_1
X_12936_ _00828_ _05995_ VPWR VGND _06033_ sg13g2_xnor2_1
X_12937_ _06021_ _06033_ VPWR VGND \atbs_core_0.n206_o[8]\ sg13g2_nor2_1
X_12938_ _00828_ _05995_ VPWR VGND _06034_ sg13g2_nand2_1
X_12939_ _00827_ _06034_ VPWR VGND _06035_ sg13g2_xor2_1
X_12940_ _06021_ _06035_ VPWR VGND \atbs_core_0.n206_o[9]\ sg13g2_nor2_1
X_12941_ _00844_ _05987_ VPWR VGND _06036_ sg13g2_nor2_1
X_12942_ _01069_ _05479_ VPWR VGND _06037_ sg13g2_nand2_1
X_12943_ _01069_ _00844_ VPWR VGND _06038_ sg13g2_nor2_1
X_12944_ _04985_ _06038_ _05475_ VPWR VGND _06039_ sg13g2_nand3_1
X_12945_ _06037_ _06039_ VPWR VGND _06040_ sg13g2_nand2_1
X_12946_ _00843_ _05475_ VPWR VGND _06041_ sg13g2_nand2_1
X_12947_ _01069_ _06041_ _06038_ VPWR VGND _06042_ sg13g2_a21o_1
X_12948_ _00846_ _06040_ _06042_ _05479_ VPWR VGND 
+ _06043_
+ sg13g2_a22oi_1
X_12949_ _01093_ _06036_ _06043_ VPWR VGND \atbs_core_0.n391_o[1]\ sg13g2_o21ai_1
X_12950_ _00846_ _04985_ _05478_ _06041_ VPWR VGND 
+ _06044_
+ sg13g2_nor4_1
X_12951_ _04985_ _00844_ _06044_ VPWR VGND _06045_ sg13g2_a21oi_1
X_12952_ _06038_ _05987_ _04985_ VPWR VGND _06046_ sg13g2_o21ai_1
X_12953_ _01071_ _06045_ _06046_ VPWR VGND \atbs_core_0.n391_o[2]\ sg13g2_o21ai_1
X_12954_ _01097_ _05282_ VPWR VGND \atbs_core_0.spike_encoder_0.n1839_o\ sg13g2_and2_1
X_12955_ _01097_ _00902_ VPWR VGND \atbs_core_0.spike_encoder_0.n1845_o\ sg13g2_and2_1
X_12956_ _00986_ VPWR VGND _06047_ sg13g2_buf_1
X_12957_ \atbs_core_0.spike_memory_0.n1953_o[0]\ \atbs_core_0.spike_memory_0.n1954_o[0]\ _06047_ VPWR VGND _06048_ sg13g2_mux2_1
X_12958_ \atbs_core_0.spike_memory_0.n1971_q[57]\ \atbs_core_0.spike_memory_0.n1953_o[0]\ _05220_ VPWR VGND _06049_ sg13g2_mux2_1
X_12959_ _00986_ VPWR VGND _06050_ sg13g2_buf_1
X_12960_ \atbs_core_0.spike_memory_0.n1955_o[0]\ \atbs_core_0.spike_memory_0.n1971_q[57]\ _06050_ VPWR VGND _06051_ sg13g2_mux2_1
X_12961_ _00986_ VPWR VGND _06052_ sg13g2_buf_1
X_12962_ \atbs_core_0.spike_memory_0.n1954_o[0]\ \atbs_core_0.spike_memory_0.n1955_o[0]\ _06052_ VPWR VGND _06053_ sg13g2_mux2_1
X_12963_ _00984_ VPWR VGND _06054_ sg13g2_buf_1
X_12964_ _06054_ VPWR VGND _06055_ sg13g2_buf_1
X_12965_ _06048_ _06049_ _06051_ _06053_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[0]\ sg13g2_mux4_1
X_12966_ \atbs_core_0.spike_memory_0.n1953_o[10]\ \atbs_core_0.spike_memory_0.n1954_o[10]\ _06047_ VPWR VGND _06056_ sg13g2_mux2_1
X_12967_ \atbs_core_0.spike_memory_0.n1971_q[67]\ \atbs_core_0.spike_memory_0.n1953_o[10]\ _05220_ VPWR VGND _06057_ sg13g2_mux2_1
X_12968_ _00986_ VPWR VGND _06058_ sg13g2_buf_1
X_12969_ \atbs_core_0.spike_memory_0.n1955_o[10]\ \atbs_core_0.spike_memory_0.n1971_q[67]\ _06058_ VPWR VGND _06059_ sg13g2_mux2_1
X_12970_ \atbs_core_0.spike_memory_0.n1954_o[10]\ \atbs_core_0.spike_memory_0.n1955_o[10]\ _06052_ VPWR VGND _06060_ sg13g2_mux2_1
X_12971_ _06056_ _06057_ _06059_ _06060_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[10]\ sg13g2_mux4_1
X_12972_ \atbs_core_0.spike_memory_0.n1953_o[11]\ \atbs_core_0.spike_memory_0.n1954_o[11]\ _06047_ VPWR VGND _06061_ sg13g2_mux2_1
X_12973_ \atbs_core_0.spike_memory_0.n1971_q[68]\ \atbs_core_0.spike_memory_0.n1953_o[11]\ _05220_ VPWR VGND _06062_ sg13g2_mux2_1
X_12974_ \atbs_core_0.spike_memory_0.n1955_o[11]\ \atbs_core_0.spike_memory_0.n1971_q[68]\ _06058_ VPWR VGND _06063_ sg13g2_mux2_1
X_12975_ \atbs_core_0.spike_memory_0.n1954_o[11]\ \atbs_core_0.spike_memory_0.n1955_o[11]\ _06052_ VPWR VGND _06064_ sg13g2_mux2_1
X_12976_ _06061_ _06062_ _06063_ _06064_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[11]\ sg13g2_mux4_1
X_12977_ \atbs_core_0.spike_memory_0.n1953_o[12]\ \atbs_core_0.spike_memory_0.n1954_o[12]\ _06047_ VPWR VGND _06065_ sg13g2_mux2_1
X_12978_ \atbs_core_0.spike_memory_0.n1971_q[69]\ \atbs_core_0.spike_memory_0.n1953_o[12]\ _05220_ VPWR VGND _06066_ sg13g2_mux2_1
X_12979_ \atbs_core_0.spike_memory_0.n1955_o[12]\ \atbs_core_0.spike_memory_0.n1971_q[69]\ _06058_ VPWR VGND _06067_ sg13g2_mux2_1
X_12980_ \atbs_core_0.spike_memory_0.n1954_o[12]\ \atbs_core_0.spike_memory_0.n1955_o[12]\ _06052_ VPWR VGND _06068_ sg13g2_mux2_1
X_12981_ _06065_ _06066_ _06067_ _06068_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[12]\ sg13g2_mux4_1
X_12982_ \atbs_core_0.spike_memory_0.n1953_o[13]\ \atbs_core_0.spike_memory_0.n1954_o[13]\ _06047_ VPWR VGND _06069_ sg13g2_mux2_1
X_12983_ \atbs_core_0.spike_memory_0.n1971_q[70]\ \atbs_core_0.spike_memory_0.n1953_o[13]\ _05220_ VPWR VGND _06070_ sg13g2_mux2_1
X_12984_ \atbs_core_0.spike_memory_0.n1955_o[13]\ \atbs_core_0.spike_memory_0.n1971_q[70]\ _06058_ VPWR VGND _06071_ sg13g2_mux2_1
X_12985_ \atbs_core_0.spike_memory_0.n1954_o[13]\ \atbs_core_0.spike_memory_0.n1955_o[13]\ _06052_ VPWR VGND _06072_ sg13g2_mux2_1
X_12986_ _06069_ _06070_ _06071_ _06072_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[13]\ sg13g2_mux4_1
X_12987_ \atbs_core_0.spike_memory_0.n1953_o[14]\ \atbs_core_0.spike_memory_0.n1954_o[14]\ _06047_ VPWR VGND _06073_ sg13g2_mux2_1
X_12988_ \atbs_core_0.spike_memory_0.n1971_q[71]\ \atbs_core_0.spike_memory_0.n1953_o[14]\ _05220_ VPWR VGND _06074_ sg13g2_mux2_1
X_12989_ \atbs_core_0.spike_memory_0.n1955_o[14]\ \atbs_core_0.spike_memory_0.n1971_q[71]\ _06058_ VPWR VGND _06075_ sg13g2_mux2_1
X_12990_ \atbs_core_0.spike_memory_0.n1954_o[14]\ \atbs_core_0.spike_memory_0.n1955_o[14]\ _06052_ VPWR VGND _06076_ sg13g2_mux2_1
X_12991_ _06073_ _06074_ _06075_ _06076_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[14]\ sg13g2_mux4_1
X_12992_ \atbs_core_0.spike_memory_0.n1953_o[15]\ \atbs_core_0.spike_memory_0.n1954_o[15]\ _06047_ VPWR VGND _06077_ sg13g2_mux2_1
X_12993_ \atbs_core_0.spike_memory_0.n1971_q[72]\ \atbs_core_0.spike_memory_0.n1953_o[15]\ _05220_ VPWR VGND _06078_ sg13g2_mux2_1
X_12994_ \atbs_core_0.spike_memory_0.n1955_o[15]\ \atbs_core_0.spike_memory_0.n1971_q[72]\ _06058_ VPWR VGND _06079_ sg13g2_mux2_1
X_12995_ \atbs_core_0.spike_memory_0.n1954_o[15]\ \atbs_core_0.spike_memory_0.n1955_o[15]\ _06052_ VPWR VGND _06080_ sg13g2_mux2_1
X_12996_ _06077_ _06078_ _06079_ _06080_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[15]\ sg13g2_mux4_1
X_12997_ \atbs_core_0.spike_memory_0.n1953_o[16]\ \atbs_core_0.spike_memory_0.n1954_o[16]\ _06047_ VPWR VGND _06081_ sg13g2_mux2_1
X_12998_ \atbs_core_0.spike_memory_0.n1971_q[73]\ \atbs_core_0.spike_memory_0.n1953_o[16]\ _05220_ VPWR VGND _06082_ sg13g2_mux2_1
X_12999_ \atbs_core_0.spike_memory_0.n1955_o[16]\ \atbs_core_0.spike_memory_0.n1971_q[73]\ _06058_ VPWR VGND _06083_ sg13g2_mux2_1
X_13000_ \atbs_core_0.spike_memory_0.n1954_o[16]\ \atbs_core_0.spike_memory_0.n1955_o[16]\ _06052_ VPWR VGND _06084_ sg13g2_mux2_1
X_13001_ _06081_ _06082_ _06083_ _06084_ _05222_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[16]\ sg13g2_mux4_1
X_13002_ \atbs_core_0.spike_memory_0.n1953_o[17]\ \atbs_core_0.spike_memory_0.n1954_o[17]\ _06047_ VPWR VGND _06085_ sg13g2_mux2_1
X_13003_ _05219_ VPWR VGND _06086_ sg13g2_buf_1
X_13004_ \atbs_core_0.spike_memory_0.n1971_q[74]\ \atbs_core_0.spike_memory_0.n1953_o[17]\ _06086_ VPWR VGND _06087_ sg13g2_mux2_1
X_13005_ \atbs_core_0.spike_memory_0.n1955_o[17]\ \atbs_core_0.spike_memory_0.n1971_q[74]\ _06058_ VPWR VGND _06088_ sg13g2_mux2_1
X_13006_ \atbs_core_0.spike_memory_0.n1954_o[17]\ \atbs_core_0.spike_memory_0.n1955_o[17]\ _06052_ VPWR VGND _06089_ sg13g2_mux2_1
X_13007_ _00985_ VPWR VGND _06090_ sg13g2_buf_1
X_13008_ _06085_ _06087_ _06088_ _06089_ _06090_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[17]\ sg13g2_mux4_1
X_13009_ _00986_ VPWR VGND _06091_ sg13g2_buf_1
X_13010_ \atbs_core_0.spike_memory_0.n1953_o[18]\ \atbs_core_0.spike_memory_0.n1954_o[18]\ _06091_ VPWR VGND _06092_ sg13g2_mux2_1
X_13011_ \atbs_core_0.spike_memory_0.n1971_q[75]\ \atbs_core_0.spike_memory_0.n1953_o[18]\ _06086_ VPWR VGND _06093_ sg13g2_mux2_1
X_13012_ \atbs_core_0.spike_memory_0.n1955_o[18]\ \atbs_core_0.spike_memory_0.n1971_q[75]\ _06058_ VPWR VGND _06094_ sg13g2_mux2_1
X_13013_ \atbs_core_0.spike_memory_0.n1954_o[18]\ \atbs_core_0.spike_memory_0.n1955_o[18]\ _06052_ VPWR VGND _06095_ sg13g2_mux2_1
X_13014_ _06092_ _06093_ _06094_ _06095_ _06090_ _06055_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[18]\ sg13g2_mux4_1
X_13015_ \atbs_core_0.spike_memory_0.n1953_o[1]\ \atbs_core_0.spike_memory_0.n1954_o[1]\ _06091_ VPWR VGND _06096_ sg13g2_mux2_1
X_13016_ \atbs_core_0.spike_memory_0.n1971_q[58]\ \atbs_core_0.spike_memory_0.n1953_o[1]\ _06086_ VPWR VGND _06097_ sg13g2_mux2_1
X_13017_ \atbs_core_0.spike_memory_0.n1955_o[1]\ \atbs_core_0.spike_memory_0.n1971_q[58]\ _06058_ VPWR VGND _06098_ sg13g2_mux2_1
X_13018_ \atbs_core_0.spike_memory_0.n1954_o[1]\ \atbs_core_0.spike_memory_0.n1955_o[1]\ _06050_ VPWR VGND _06099_ sg13g2_mux2_1
X_13019_ _06096_ _06097_ _06098_ _06099_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[1]\ sg13g2_mux4_1
X_13020_ \atbs_core_0.spike_memory_0.n1953_o[2]\ \atbs_core_0.spike_memory_0.n1954_o[2]\ _06091_ VPWR VGND _06100_ sg13g2_mux2_1
X_13021_ \atbs_core_0.spike_memory_0.n1971_q[59]\ \atbs_core_0.spike_memory_0.n1953_o[2]\ _06086_ VPWR VGND _06101_ sg13g2_mux2_1
X_13022_ \atbs_core_0.spike_memory_0.n1955_o[2]\ \atbs_core_0.spike_memory_0.n1971_q[59]\ _05219_ VPWR VGND _06102_ sg13g2_mux2_1
X_13023_ \atbs_core_0.spike_memory_0.n1954_o[2]\ \atbs_core_0.spike_memory_0.n1955_o[2]\ _06050_ VPWR VGND _06103_ sg13g2_mux2_1
X_13024_ _06100_ _06101_ _06102_ _06103_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[2]\ sg13g2_mux4_1
X_13025_ \atbs_core_0.spike_memory_0.n1953_o[3]\ \atbs_core_0.spike_memory_0.n1954_o[3]\ _06091_ VPWR VGND _06104_ sg13g2_mux2_1
X_13026_ \atbs_core_0.spike_memory_0.n1971_q[60]\ \atbs_core_0.spike_memory_0.n1953_o[3]\ _06086_ VPWR VGND _06105_ sg13g2_mux2_1
X_13027_ \atbs_core_0.spike_memory_0.n1955_o[3]\ \atbs_core_0.spike_memory_0.n1971_q[60]\ _05219_ VPWR VGND _06106_ sg13g2_mux2_1
X_13028_ \atbs_core_0.spike_memory_0.n1954_o[3]\ \atbs_core_0.spike_memory_0.n1955_o[3]\ _06050_ VPWR VGND _06107_ sg13g2_mux2_1
X_13029_ _06104_ _06105_ _06106_ _06107_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[3]\ sg13g2_mux4_1
X_13030_ \atbs_core_0.spike_memory_0.n1953_o[4]\ \atbs_core_0.spike_memory_0.n1954_o[4]\ _06091_ VPWR VGND _06108_ sg13g2_mux2_1
X_13031_ \atbs_core_0.spike_memory_0.n1971_q[61]\ \atbs_core_0.spike_memory_0.n1953_o[4]\ _06086_ VPWR VGND _06109_ sg13g2_mux2_1
X_13032_ \atbs_core_0.spike_memory_0.n1955_o[4]\ \atbs_core_0.spike_memory_0.n1971_q[61]\ _05219_ VPWR VGND _06110_ sg13g2_mux2_1
X_13033_ \atbs_core_0.spike_memory_0.n1954_o[4]\ \atbs_core_0.spike_memory_0.n1955_o[4]\ _06050_ VPWR VGND _06111_ sg13g2_mux2_1
X_13034_ _06108_ _06109_ _06110_ _06111_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[4]\ sg13g2_mux4_1
X_13035_ \atbs_core_0.spike_memory_0.n1953_o[5]\ \atbs_core_0.spike_memory_0.n1954_o[5]\ _06091_ VPWR VGND _06112_ sg13g2_mux2_1
X_13036_ \atbs_core_0.spike_memory_0.n1971_q[62]\ \atbs_core_0.spike_memory_0.n1953_o[5]\ _06086_ VPWR VGND _06113_ sg13g2_mux2_1
X_13037_ \atbs_core_0.spike_memory_0.n1955_o[5]\ \atbs_core_0.spike_memory_0.n1971_q[62]\ _05219_ VPWR VGND _06114_ sg13g2_mux2_1
X_13038_ \atbs_core_0.spike_memory_0.n1954_o[5]\ \atbs_core_0.spike_memory_0.n1955_o[5]\ _06050_ VPWR VGND _06115_ sg13g2_mux2_1
X_13039_ _06112_ _06113_ _06114_ _06115_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[5]\ sg13g2_mux4_1
X_13040_ \atbs_core_0.spike_memory_0.n1953_o[6]\ \atbs_core_0.spike_memory_0.n1954_o[6]\ _06091_ VPWR VGND _06116_ sg13g2_mux2_1
X_13041_ \atbs_core_0.spike_memory_0.n1971_q[63]\ \atbs_core_0.spike_memory_0.n1953_o[6]\ _06086_ VPWR VGND _06117_ sg13g2_mux2_1
X_13042_ \atbs_core_0.spike_memory_0.n1955_o[6]\ \atbs_core_0.spike_memory_0.n1971_q[63]\ _05219_ VPWR VGND _06118_ sg13g2_mux2_1
X_13043_ \atbs_core_0.spike_memory_0.n1954_o[6]\ \atbs_core_0.spike_memory_0.n1955_o[6]\ _06050_ VPWR VGND _06119_ sg13g2_mux2_1
X_13044_ _06116_ _06117_ _06118_ _06119_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[6]\ sg13g2_mux4_1
X_13045_ \atbs_core_0.spike_memory_0.n1953_o[7]\ \atbs_core_0.spike_memory_0.n1954_o[7]\ _06091_ VPWR VGND _06120_ sg13g2_mux2_1
X_13046_ \atbs_core_0.spike_memory_0.n1971_q[64]\ \atbs_core_0.spike_memory_0.n1953_o[7]\ _06086_ VPWR VGND _06121_ sg13g2_mux2_1
X_13047_ \atbs_core_0.spike_memory_0.n1955_o[7]\ \atbs_core_0.spike_memory_0.n1971_q[64]\ _05219_ VPWR VGND _06122_ sg13g2_mux2_1
X_13048_ \atbs_core_0.spike_memory_0.n1954_o[7]\ \atbs_core_0.spike_memory_0.n1955_o[7]\ _06050_ VPWR VGND _06123_ sg13g2_mux2_1
X_13049_ _06120_ _06121_ _06122_ _06123_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[7]\ sg13g2_mux4_1
X_13050_ \atbs_core_0.spike_memory_0.n1953_o[8]\ \atbs_core_0.spike_memory_0.n1954_o[8]\ _06091_ VPWR VGND _06124_ sg13g2_mux2_1
X_13051_ \atbs_core_0.spike_memory_0.n1971_q[65]\ \atbs_core_0.spike_memory_0.n1953_o[8]\ _06086_ VPWR VGND _06125_ sg13g2_mux2_1
X_13052_ \atbs_core_0.spike_memory_0.n1955_o[8]\ \atbs_core_0.spike_memory_0.n1971_q[65]\ _05219_ VPWR VGND _06126_ sg13g2_mux2_1
X_13053_ \atbs_core_0.spike_memory_0.n1954_o[8]\ \atbs_core_0.spike_memory_0.n1955_o[8]\ _06050_ VPWR VGND _06127_ sg13g2_mux2_1
X_13054_ _06124_ _06125_ _06126_ _06127_ _06090_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[8]\ sg13g2_mux4_1
X_13055_ \atbs_core_0.spike_memory_0.n1953_o[9]\ \atbs_core_0.spike_memory_0.n1954_o[9]\ _06091_ VPWR VGND _06128_ sg13g2_mux2_1
X_13056_ \atbs_core_0.spike_memory_0.n1971_q[66]\ \atbs_core_0.spike_memory_0.n1953_o[9]\ _06047_ VPWR VGND _06129_ sg13g2_mux2_1
X_13057_ \atbs_core_0.spike_memory_0.n1955_o[9]\ \atbs_core_0.spike_memory_0.n1971_q[66]\ _05219_ VPWR VGND _06130_ sg13g2_mux2_1
X_13058_ \atbs_core_0.spike_memory_0.n1954_o[9]\ \atbs_core_0.spike_memory_0.n1955_o[9]\ _06050_ VPWR VGND _06131_ sg13g2_mux2_1
X_13059_ _06128_ _06129_ _06130_ _06131_ _00985_ _06054_ 
+ VPWR
+ VGND \atbs_core_0.spike_memory_0.n1985_o[9]\ sg13g2_mux4_1
X_13060_ _01795_ _01970_ _01788_ VPWR VGND _06132_ sg13g2_nand3_1
X_13061_ _02222_ _06132_ VPWR VGND _06133_ sg13g2_nor2_1
X_13062_ _01810_ _01784_ _06133_ VPWR VGND _06134_ sg13g2_nand3_1
X_13063_ _01983_ _06134_ VPWR VGND _06135_ sg13g2_or2_1
X_13064_ _05194_ _06135_ VPWR VGND _06136_ sg13g2_nor2_1
X_13065_ _01998_ _05100_ _06136_ VPWR VGND _06137_ sg13g2_nand3_1
X_13066_ _01728_ _06137_ VPWR VGND _06138_ sg13g2_nor2_1
X_13067_ _01954_ _05117_ _06138_ VPWR VGND _06139_ sg13g2_nand3_1
X_13068_ _05134_ _06139_ VPWR VGND _06140_ sg13g2_nor2_1
X_13069_ _02049_ _05147_ _06140_ VPWR VGND _06141_ sg13g2_nand3_1
X_13070_ _01895_ _03396_ _06141_ VPWR VGND \atbs_core_0.time_measurement_0.n1809_o\ sg13g2_nor3_1
X_13071_ _05118_ \atbs_core_0.time_measurement_0.n1809_o\ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[0]\ sg13g2_nor2_1
X_13072_ _02250_ _06137_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[10]\ sg13g2_xnor2_1
X_13073_ _05117_ _06138_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[11]\ sg13g2_xor2_1
X_13074_ _05117_ _06138_ VPWR VGND _06142_ sg13g2_nand2_1
X_13075_ _01954_ _06142_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[12]\ sg13g2_xnor2_1
X_13076_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[13]\ _06139_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[13]\ sg13g2_xnor2_1
X_13077_ _01703_ _06140_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[14]\ sg13g2_xnor2_1
X_13078_ _02049_ _06140_ VPWR VGND _06143_ sg13g2_nand2_1
X_13079_ _05147_ _06143_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[15]\ sg13g2_xnor2_1
X_13080_ _02069_ _06141_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[16]\ sg13g2_xnor2_1
X_13081_ _03396_ _06141_ VPWR VGND _06144_ sg13g2_nor2_1
X_13082_ _01895_ _06144_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[17]\ sg13g2_xnor2_1
X_13083_ _01795_ _01970_ VPWR VGND _06145_ sg13g2_nand2_1
X_13084_ _02382_ _06145_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[2]\ sg13g2_xnor2_1
X_13085_ _01803_ _06132_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[3]\ sg13g2_xnor2_1
X_13086_ _01964_ _06133_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[4]\ sg13g2_xnor2_1
X_13087_ _01784_ _06133_ VPWR VGND _06146_ sg13g2_nand2_1
X_13088_ _01810_ _06146_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[5]\ sg13g2_xnor2_1
X_13089_ _01827_ _06134_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[6]\ sg13g2_xnor2_1
X_13090_ _05102_ _06135_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[7]\ sg13g2_xnor2_1
X_13091_ _04239_ _06136_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[8]\ sg13g2_xnor2_1
X_13092_ _01998_ _06136_ VPWR VGND _06147_ sg13g2_nand2_1
X_13093_ _05100_ _06147_ VPWR VGND \atbs_core_0.time_measurement_0.n1813_o[9]\ sg13g2_xnor2_1
X_13094_ _00758_ VPWR VGND _06148_ sg13g2_inv_1
X_13095_ _00759_ VPWR VGND _06149_ sg13g2_inv_1
X_13096_ _00773_ _00774_ VPWR VGND _06150_ sg13g2_nand2b_1
X_13097_ _00771_ _06150_ VPWR VGND _06151_ sg13g2_nand2_1
X_13098_ _00767_ _06151_ VPWR VGND _06152_ sg13g2_nand2_1
X_13099_ _00771_ _06150_ _06152_ VPWR VGND _06153_ sg13g2_o21ai_1
X_13100_ _00750_ _00766_ _06153_ VPWR VGND _06154_ sg13g2_o21ai_1
X_13101_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ VPWR VGND _06155_ sg13g2_inv_1
X_13102_ _00767_ _06155_ _00764_ VPWR VGND _06156_ sg13g2_o21ai_1
X_13103_ _00770_ _06154_ _06156_ _00765_ VPWR VGND 
+ _06157_
+ sg13g2_a22oi_1
X_13104_ _06157_ _00755_ VPWR VGND _06158_ sg13g2_nand2b_1
X_13105_ _00755_ _06157_ VPWR VGND _06159_ sg13g2_nor2b_1
X_13106_ _00758_ _06149_ _06158_ _00754_ _06159_ VPWR 
+ VGND
+ _06160_ sg13g2_a221oi_1
X_13107_ _06148_ _00759_ _00780_ _00777_ _06160_ VPWR 
+ VGND
+ _06161_ sg13g2_a221oi_1
X_13108_ _00754_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ VPWR VGND _06162_ sg13g2_nand2b_1
X_13109_ _00781_ _06161_ _06162_ VPWR VGND _06163_ sg13g2_o21ai_1
X_13110_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ _00754_ VPWR VGND _06164_ sg13g2_nand2b_1
X_13111_ _06163_ _06164_ _00971_ VPWR VGND _06165_ sg13g2_a21o_1
X_13112_ _06165_ VPWR VGND _06166_ sg13g2_buf_1
X_13113_ _00773_ _06166_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[0]\ sg13g2_nor2_1
X_13114_ _00773_ _00771_ VPWR VGND _06167_ sg13g2_xnor2_1
X_13115_ _06166_ _06167_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[1]\ sg13g2_nor2_1
X_13116_ _00773_ _00771_ VPWR VGND _06168_ sg13g2_nand2_1
X_13117_ _00766_ _06168_ VPWR VGND _06169_ sg13g2_xnor2_1
X_13118_ _06166_ _06169_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[2]\ sg13g2_nor2_1
X_13119_ _00773_ _00771_ _00752_ VPWR VGND _06170_ sg13g2_nand3_1
X_13120_ _06155_ _06170_ VPWR VGND _06171_ sg13g2_xnor2_1
X_13121_ _06166_ _06171_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[3]\ sg13g2_nor2_1
X_13122_ _06155_ _06170_ VPWR VGND _06172_ sg13g2_nor2_1
X_13123_ _00763_ _06172_ VPWR VGND _06173_ sg13g2_xnor2_1
X_13124_ _06166_ _06173_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[4]\ sg13g2_nor2_1
X_13125_ _00763_ _06172_ VPWR VGND _06174_ sg13g2_nand2_1
X_13126_ _00755_ _06174_ VPWR VGND _06175_ sg13g2_xor2_1
X_13127_ _06166_ _06175_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[5]\ sg13g2_nor2_1
X_13128_ _00763_ _00755_ _06172_ VPWR VGND _06176_ sg13g2_nand3_1
X_13129_ _06149_ _06176_ VPWR VGND _06177_ sg13g2_xnor2_1
X_13130_ _06166_ _06177_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[6]\ sg13g2_nor2_1
X_13131_ _06149_ _06176_ VPWR VGND _06178_ sg13g2_or2_1
X_13132_ _00778_ _06178_ VPWR VGND _06179_ sg13g2_xnor2_1
X_13133_ _06166_ _06179_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[7]\ sg13g2_nor2_1
X_13134_ _00778_ _06178_ VPWR VGND _06180_ sg13g2_nor2_1
X_13135_ _00006_ _06180_ VPWR VGND _06181_ sg13g2_xnor2_1
X_13136_ _06166_ _06181_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n2836_o[8]\ sg13g2_nor2b_1
X_13137_ _00956_ _05489_ VPWR VGND _06182_ sg13g2_nand2_1
X_13138_ _00748_ _00971_ _00789_ _06182_ VPWR VGND 
+ \atbs_core_0.uart_0.uart_rx_0.n2880_o\
+ sg13g2_nor4_1
X_13139_ _00754_ _00798_ VPWR VGND _06183_ sg13g2_nand2b_1
X_13140_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ VPWR VGND _06184_ sg13g2_inv_1
X_13141_ _00797_ _00754_ VPWR VGND _06185_ sg13g2_nand2b_1
X_13142_ _00774_ VPWR VGND _06186_ sg13g2_inv_1
X_13143_ _06186_ _00809_ _00801_ VPWR VGND _06187_ sg13g2_o21ai_1
X_13144_ _06186_ _00809_ _00801_ _00802_ VPWR VGND 
+ _06188_
+ sg13g2_nor4_1
X_13145_ _00767_ _06187_ _06188_ VPWR VGND _06189_ sg13g2_a21o_1
X_13146_ _00802_ _00807_ VPWR VGND _06190_ sg13g2_nand2_1
X_13147_ \atbs_core_0.baudrate_adj_uart[1]\ _06190_ VPWR VGND _06191_ sg13g2_nand2_1
X_13148_ _00802_ _00807_ _06191_ VPWR VGND _06192_ sg13g2_o21ai_1
X_13149_ _00806_ _06189_ _06192_ VPWR VGND _06193_ sg13g2_a21o_1
X_13150_ _00795_ _06193_ VPWR VGND _06194_ sg13g2_nor2b_1
X_13151_ _06193_ _00795_ VPWR VGND _06195_ sg13g2_nand2b_1
X_13152_ _00762_ _06194_ _06195_ VPWR VGND _06196_ sg13g2_o21ai_1
X_13153_ _00754_ _00797_ VPWR VGND _06197_ sg13g2_nor2b_1
X_13154_ _06148_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ _06185_ _06196_ _06197_ VPWR 
+ VGND
+ _06198_ sg13g2_a221oi_1
X_13155_ _00758_ _06184_ _06198_ VPWR VGND _06199_ sg13g2_a21oi_1
X_13156_ _00793_ _06199_ _00780_ VPWR VGND _06200_ sg13g2_a21o_1
X_13157_ _00793_ _06199_ _06200_ VPWR VGND _06201_ sg13g2_o21ai_1
X_13158_ _00798_ _00754_ VPWR VGND _06202_ sg13g2_nor2b_1
X_13159_ _06183_ _06201_ _06202_ VPWR VGND _06203_ sg13g2_a21oi_1
X_13160_ _06203_ VPWR VGND _06204_ sg13g2_buf_1
X_13161_ _00809_ _06204_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[0]\ sg13g2_nor2_1
X_13162_ _00809_ _00801_ VPWR VGND _06205_ sg13g2_xnor2_1
X_13163_ _06204_ _06205_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[1]\ sg13g2_nor2_1
X_13164_ _00809_ _00801_ VPWR VGND _06206_ sg13g2_nand2_1
X_13165_ _00805_ _06206_ VPWR VGND _06207_ sg13g2_xor2_1
X_13166_ _06204_ _06207_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[2]\ sg13g2_nor2_1
X_13167_ _00802_ VPWR VGND _06208_ sg13g2_inv_1
X_13168_ _00809_ _00801_ _00805_ VPWR VGND _06209_ sg13g2_nand3_1
X_13169_ _06208_ _06209_ VPWR VGND _06210_ sg13g2_xnor2_1
X_13170_ _06204_ _06210_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[3]\ sg13g2_nor2_1
X_13171_ _06208_ _06209_ VPWR VGND _06211_ sg13g2_nor2_1
X_13172_ _00795_ _06211_ VPWR VGND _06212_ sg13g2_xnor2_1
X_13173_ _06204_ _06212_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[4]\ sg13g2_nor2_1
X_13174_ _00795_ _06211_ VPWR VGND _06213_ sg13g2_nand2_1
X_13175_ _00797_ _06213_ VPWR VGND _06214_ sg13g2_xor2_1
X_13176_ _06204_ _06214_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[5]\ sg13g2_nor2_1
X_13177_ _00797_ _00795_ _06211_ VPWR VGND _06215_ sg13g2_nand3_1
X_13178_ _06184_ _06215_ VPWR VGND _06216_ sg13g2_xnor2_1
X_13179_ _06204_ _06216_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[6]\ sg13g2_nor2_1
X_13180_ _00793_ VPWR VGND _06217_ sg13g2_inv_1
X_13181_ _06184_ _06215_ VPWR VGND _06218_ sg13g2_or2_1
X_13182_ _06217_ _06218_ VPWR VGND _06219_ sg13g2_xnor2_1
X_13183_ _06204_ _06219_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[7]\ sg13g2_nor2_1
X_13184_ _06217_ _06218_ VPWR VGND _06220_ sg13g2_nor2_1
X_13185_ _00798_ _06220_ VPWR VGND _06221_ sg13g2_xnor2_1
X_13186_ _06204_ _06221_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n2712_o[8]\ sg13g2_nor2_1
X_13187_ _00817_ _00978_ _00791_ _00815_ VPWR VGND 
+ \atbs_core_0.uart_0.uart_tx_0.n2776_o\
+ sg13g2_nor4_1
X_13188_ _00974_ _00975_ VPWR VGND _06222_ sg13g2_nor2_1
X_13189_ \atbs_core_0.uart_0.uart_tx_0.n2787_o\ _00976_ VPWR VGND _06223_ sg13g2_nand2b_1
X_13190_ _00976_ \atbs_core_0.uart_0.uart_tx_0.n2783_o\ _06223_ VPWR VGND _06224_ sg13g2_o21ai_1
X_13191_ _00816_ _00791_ VPWR VGND _06225_ sg13g2_xor2_1
X_13192_ _00022_ VPWR VGND _06226_ sg13g2_inv_1
X_13193_ \atbs_core_0.uart_0.uart_tx_0.n2721_o\ _00978_ _06226_ VPWR VGND _06227_ sg13g2_nor3_1
X_13194_ _06222_ _06224_ _06225_ _06227_ VPWR VGND 
+ _06228_
+ sg13g2_a22oi_1
X_13195_ _00974_ \atbs_core_0.uart_0.uart_tx_0.n2786_o\ VPWR VGND _06229_ sg13g2_nand2_1
X_13196_ _00974_ \atbs_core_0.uart_0.uart_tx_0.n2784_o\ VPWR VGND _06230_ sg13g2_nand2b_1
X_13197_ _00975_ _06229_ _06230_ VPWR VGND _06231_ sg13g2_nand3_1
X_13198_ _00975_ \atbs_core_0.uart_0.uart_tx_0.n2785_o\ _06231_ VPWR VGND _06232_ sg13g2_o21ai_1
X_13199_ \atbs_core_0.uart_0.uart_tx_0.n2789_o\ VPWR VGND _06233_ sg13g2_inv_1
X_13200_ _00974_ _00975_ \atbs_core_0.uart_0.uart_tx_0.n2790_o\ VPWR VGND _06234_ sg13g2_nand3_1
X_13201_ _00975_ _06233_ _06234_ VPWR VGND _06235_ sg13g2_o21ai_1
X_13202_ _00976_ \atbs_core_0.uart_0.uart_tx_0.n2788_o\ VPWR VGND _06236_ sg13g2_nand2_1
X_13203_ _00975_ _06236_ _00974_ VPWR VGND _06237_ sg13g2_a21oi_1
X_13204_ _00976_ _06235_ _06237_ VPWR VGND _06238_ sg13g2_a21oi_1
X_13205_ _00976_ _06232_ _06238_ VPWR VGND _06239_ sg13g2_o21ai_1
X_13206_ _00816_ _00022_ _00814_ VPWR VGND _06240_ sg13g2_nand3_1
X_13207_ _00817_ _00816_ _06240_ VPWR VGND _06241_ sg13g2_o21ai_1
X_13208_ \atbs_core_0.uart_0.uart_tx_0.n2758_o\ _00818_ _00816_ VPWR VGND _06242_ sg13g2_nor3_1
X_13209_ _00818_ _06241_ _06242_ VPWR VGND _06243_ sg13g2_a21oi_1
X_13210_ _00978_ _00791_ _06243_ VPWR VGND _06244_ sg13g2_nor3_1
X_13211_ _06228_ _06239_ _06244_ VPWR VGND uart_tx_o sg13g2_a21o_1
X_13212_ _06940_ VPWR VGND sg13g2_tiehi
X\atbs_core_0.adaptive_ctrl_0.n1441_q$_DFFE_PP0P_  clock_i _00125_ \atbs_core_0.adaptive_ctrl_0.adapt_on_overflow\ _00029_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1442_q$_DFFE_PP0P_  clock_i _00126_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _06934_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1443_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1345_o\ \atbs_core_0.adaptive_ctrl_0.adaptive_strb\ _00024_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1444_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1348_o\ \atbs_core_0.adaptive_ctrl_0.n1444_q\ _00023_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1445_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1352_o\ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ _06933_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[0]$_DFFE_PP1P_  clock_i _00127_ _00090_ \atbs_core_0.adaptive_ctrl_0.delta_steps[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[1]$_DFFE_PP0P_  clock_i _00128_ \atbs_core_0.adaptive_ctrl_0.delta_steps[1]\ _00045_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[2]$_DFFE_PP0P_  clock_i _00129_ \atbs_core_0.adaptive_ctrl_0.delta_steps[2]\ _00043_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[3]$_DFFE_PP0P_  clock_i _00130_ \atbs_core_0.adaptive_ctrl_0.delta_steps[3]\ _00040_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[4]$_DFFE_PP0P_  clock_i _00131_ \atbs_core_0.adaptive_ctrl_0.delta_steps[4]\ _00039_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[5]$_DFFE_PP0P_  clock_i _00132_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ _00036_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[6]$_DFFE_PP0P_  clock_i _00133_ \atbs_core_0.adaptive_ctrl_0.delta_steps[6]\ _00035_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1446_q[7]$_DFFE_PP0P_  clock_i _00134_ \atbs_core_0.adaptive_ctrl_0.delta_steps[7]\ _00032_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[0]$_DFFE_PP1P_  clock_i _00135_ _00091_ \atbs_core_0.adaptive_ctrl_0.n1447_q[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[1]$_DFFE_PP0P_  clock_i _00136_ \atbs_core_0.adaptive_ctrl_0.n1447_q[1]\ _06932_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[2]$_DFFE_PP0P_  clock_i _00137_ \atbs_core_0.adaptive_ctrl_0.n1447_q[2]\ _06931_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[3]$_DFFE_PP0P_  clock_i _00138_ \atbs_core_0.adaptive_ctrl_0.n1447_q[3]\ _06930_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[4]$_DFFE_PP0P_  clock_i _00139_ \atbs_core_0.adaptive_ctrl_0.n1447_q[4]\ _06929_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[5]$_DFFE_PP0P_  clock_i _00140_ \atbs_core_0.adaptive_ctrl_0.n1447_q[5]\ _06928_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[6]$_DFFE_PP0P_  clock_i _00141_ \atbs_core_0.adaptive_ctrl_0.n1447_q[6]\ _06927_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1447_q[7]$_DFFE_PP0P_  clock_i _00142_ \atbs_core_0.adaptive_ctrl_0.n1447_q[7]\ _06926_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[0]$_DFFE_PP1P_  clock_i _00143_ _00092_ \atbs_core_0.adaptive_ctrl_0.n1368_o[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[1]$_DFFE_PP0P_  clock_i _00144_ \atbs_core_0.adaptive_ctrl_0.n1368_o[1]\ _00046_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[2]$_DFFE_PP1P_  clock_i _00145_ _00093_ \atbs_core_0.adaptive_ctrl_0.n1368_o[2]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[3]$_DFFE_PP1P_  clock_i _00146_ _00094_ \atbs_core_0.adaptive_ctrl_0.n1368_o[3]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[4]$_DFFE_PP1P_  clock_i _00147_ _00095_ \atbs_core_0.adaptive_ctrl_0.n1368_o[4]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[5]$_DFFE_PP1P_  clock_i _00148_ _00096_ \atbs_core_0.adaptive_ctrl_0.n1368_o[5]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[6]$_DFFE_PP1P_  clock_i _00149_ _00097_ \atbs_core_0.adaptive_ctrl_0.n1368_o[6]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[7]$_DFFE_PP0P_  clock_i _00150_ \atbs_core_0.adaptive_ctrl_0.n1368_o[7]\ _00033_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1448_q[8]$_DFFE_PP0P_  clock_i _00151_ \atbs_core_0.adaptive_ctrl_0.n1448_q[8]\ _00026_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[0]$_DFFE_PP1P_  clock_i _00152_ _00098_ \atbs_core_0.adaptive_ctrl_0.n1373_o[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[1]$_DFFE_PP1P_  clock_i _00153_ _00099_ \atbs_core_0.adaptive_ctrl_0.n1373_o[1]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[2]$_DFFE_PP1P_  clock_i _00154_ _00100_ \atbs_core_0.adaptive_ctrl_0.n1373_o[2]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[3]$_DFFE_PP1P_  clock_i _00155_ _00101_ \atbs_core_0.adaptive_ctrl_0.n1373_o[3]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[4]$_DFFE_PP1P_  clock_i _00156_ _00102_ \atbs_core_0.adaptive_ctrl_0.n1373_o[4]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[5]$_DFFE_PP1P_  clock_i _00157_ _00103_ \atbs_core_0.adaptive_ctrl_0.n1373_o[5]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[6]$_DFFE_PP1P_  clock_i _00158_ _00104_ \atbs_core_0.adaptive_ctrl_0.n1373_o[6]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[7]$_DFFE_PP0P_  clock_i _00159_ \atbs_core_0.adaptive_ctrl_0.n1373_o[7]\ _00034_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1449_q[8]$_DFFE_PP0P_  clock_i _00160_ \atbs_core_0.adaptive_ctrl_0.n1449_q[8]\ _06925_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[0]$_DFFE_PP0N_  clock_i _00161_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ _06924_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[100]$_DFFE_PP0N_  clock_i _00162_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[10]\ _06923_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[101]$_DFFE_PP0N_  clock_i _00163_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[11]\ _06922_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[102]$_DFFE_PP0N_  clock_i _00164_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[12]\ _06921_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[103]$_DFFE_PP0N_  clock_i _00165_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[13]\ _06920_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[104]$_DFFE_PP0N_  clock_i _00166_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[14]\ _06919_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[105]$_DFFE_PP0N_  clock_i _00167_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[15]\ _06918_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[106]$_DFFE_PP0N_  clock_i _00168_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[16]\ _06917_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[107]$_DFFE_PP0N_  clock_i _00169_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[17]\ _06916_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[108]$_DFFE_PP0N_  clock_i _00170_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ _06915_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[109]$_DFFE_PP0N_  clock_i _00171_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[115]\ _06914_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[10]$_DFFE_PP0N_  clock_i _00172_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[10]\ _06913_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[110]$_DFFE_PP0N_  clock_i _00173_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _06912_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[111]$_DFFE_PP0N_  clock_i _00174_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ _06911_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[112]$_DFFE_PP0N_  clock_i _00175_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ _06910_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[113]$_DFFE_PP0N_  clock_i _00176_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[119]\ _06909_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[114]$_DFFE_PP0N_  clock_i _00177_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[6]\ _06908_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[115]$_DFFE_PP0N_  clock_i _00178_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[7]\ _06907_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[116]$_DFFE_PP0N_  clock_i _00179_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[8]\ _06906_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[117]$_DFFE_PP0N_  clock_i _00180_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[9]\ _06905_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[118]$_DFFE_PP0N_  clock_i _00181_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[10]\ _06904_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[119]$_DFFE_PP0N_  clock_i _00182_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[11]\ _06903_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[11]$_DFFE_PP0N_  clock_i _00183_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[11]\ _06902_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[120]$_DFFE_PP0N_  clock_i _00184_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[12]\ _06901_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[121]$_DFFE_PP0N_  clock_i _00185_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[13]\ _06900_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[122]$_DFFE_PP0N_  clock_i _00186_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[14]\ _06899_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[123]$_DFFE_PP0N_  clock_i _00187_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[15]\ _06898_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[124]$_DFFE_PP0N_  clock_i _00188_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[16]\ _06897_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[125]$_DFFE_PP0N_  clock_i _00189_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2089_o[17]\ _06896_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[126]$_DFFE_PP0N_  clock_i _00190_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ _06895_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[127]$_DFFE_PP0N_  clock_i _00191_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ _06894_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[128]$_DFFE_PP0N_  clock_i _00192_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ _06893_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[129]$_DFFE_PP0N_  clock_i _00193_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ _06892_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[12]$_DFFE_PP0N_  clock_i _00194_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[12]\ _06891_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[130]$_DFFE_PP0N_  clock_i _00195_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ _06890_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[131]$_DFFE_PP0N_  clock_i _00196_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[138]\ _06889_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[132]$_DFFE_PP0N_  clock_i _00197_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[6]\ _06888_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[133]$_DFFE_PP0N_  clock_i _00198_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[7]\ _06887_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[134]$_DFFE_PP0N_  clock_i _00199_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[8]\ _06886_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[135]$_DFFE_PP0N_  clock_i _00200_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[9]\ _06885_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[136]$_DFFE_PP0N_  clock_i _00201_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[10]\ _06884_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[137]$_DFFE_PP0N_  clock_i _00202_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[11]\ _06883_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[138]$_DFFE_PP0N_  clock_i _00203_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[12]\ _06882_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[139]$_DFFE_PP0N_  clock_i _00204_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[13]\ _06881_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[13]$_DFFE_PP0N_  clock_i _00205_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[13]\ _06880_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[140]$_DFFE_PP0N_  clock_i _00206_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[14]\ _06879_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[141]$_DFFE_PP0N_  clock_i _00207_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[15]\ _06878_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[142]$_DFFE_PP0N_  clock_i _00208_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[16]\ _06877_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[143]$_DFFE_PP0N_  clock_i _00209_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2092_o[17]\ _06876_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[144]$_DFFE_PP0N_  clock_i _00210_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ _06875_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[145]$_DFFE_PP0N_  clock_i _00211_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _06874_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[146]$_DFFE_PP0N_  clock_i _00212_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[154]\ _06873_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[147]$_DFFE_PP0N_  clock_i _00213_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ _06872_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[148]$_DFFE_PP0N_  clock_i _00214_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ _06871_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[149]$_DFFE_PP0N_  clock_i _00215_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[157]\ _06870_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[14]$_DFFE_PP0N_  clock_i _00216_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[14]\ _06869_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[150]$_DFFE_PP0N_  clock_i _00217_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[6]\ _06868_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[151]$_DFFE_PP0N_  clock_i _00218_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[7]\ _06867_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[152]$_DFFE_PP0N_  clock_i _00219_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[8]\ _06866_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[153]$_DFFE_PP0N_  clock_i _00220_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[9]\ _06865_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[154]$_DFFE_PP0N_  clock_i _00221_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[10]\ _06864_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[155]$_DFFE_PP0N_  clock_i _00222_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[11]\ _06863_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[156]$_DFFE_PP0N_  clock_i _00223_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[12]\ _06862_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[157]$_DFFE_PP0N_  clock_i _00224_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[13]\ _06861_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[158]$_DFFE_PP0N_  clock_i _00225_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[14]\ _06860_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[159]$_DFFE_PP0N_  clock_i _00226_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[15]\ _06859_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[15]$_DFFE_PP0N_  clock_i _00227_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[15]\ _06858_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[160]$_DFFE_PP0N_  clock_i _00228_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[16]\ _06857_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[161]$_DFFE_PP0N_  clock_i _00229_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2095_o[17]\ _06856_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[162]$_DFFE_PP0N_  clock_i _00230_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ _06855_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[163]$_DFFE_PP0N_  clock_i _00231_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[172]\ _06854_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[164]$_DFFE_PP0N_  clock_i _00232_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _06853_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[165]$_DFFE_PP0N_  clock_i _00233_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _06852_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[166]$_DFFE_PP0N_  clock_i _00234_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ _06851_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[167]$_DFFE_PP0N_  clock_i _00235_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[176]\ _06850_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[168]$_DFFE_PP0N_  clock_i _00236_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[6]\ _06849_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[169]$_DFFE_PP0N_  clock_i _00237_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[7]\ _06848_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[16]$_DFFE_PP0N_  clock_i _00238_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[16]\ _06847_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[170]$_DFFE_PP0N_  clock_i _00239_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[8]\ _06846_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[171]$_DFFE_PP0N_  clock_i _00240_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[9]\ _06845_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[172]$_DFFE_PP0N_  clock_i _00241_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[10]\ _06844_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[173]$_DFFE_PP0N_  clock_i _00242_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[11]\ _06843_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[174]$_DFFE_PP0N_  clock_i _00243_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[12]\ _06842_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[175]$_DFFE_PP0N_  clock_i _00244_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[13]\ _06841_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[176]$_DFFE_PP0N_  clock_i _00245_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[14]\ _06840_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[177]$_DFFE_PP0N_  clock_i _00246_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[15]\ _06839_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[178]$_DFFE_PP0N_  clock_i _00247_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[16]\ _06838_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[179]$_DFFE_PP0N_  clock_i _00248_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2098_o[17]\ _06837_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[17]$_DFFE_PP0N_  clock_i _00249_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[17]\ _06836_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[180]$_DFFE_PP0N_  clock_i _00250_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ _06835_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[181]$_DFFE_PP0N_  clock_i _00251_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[191]\ _06834_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[182]$_DFFE_PP0N_  clock_i _00252_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ _06833_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[183]$_DFFE_PP0N_  clock_i _00253_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[193]\ _06832_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[184]$_DFFE_PP0N_  clock_i _00254_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ _06831_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[185]$_DFFE_PP0N_  clock_i _00255_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ _06830_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[186]$_DFFE_PP0N_  clock_i _00256_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[6]\ _06829_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[187]$_DFFE_PP0N_  clock_i _00257_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[7]\ _06828_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[188]$_DFFE_PP0N_  clock_i _00258_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[8]\ _06827_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[189]$_DFFE_PP0N_  clock_i _00259_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[9]\ _06826_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[18]$_DFFE_PP0N_  clock_i _00260_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ _06825_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[190]$_DFFE_PP0N_  clock_i _00261_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[10]\ _06824_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[191]$_DFFE_PP0N_  clock_i _00262_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[11]\ _06823_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[192]$_DFFE_PP0N_  clock_i _00263_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[12]\ _06822_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[193]$_DFFE_PP0N_  clock_i _00264_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[13]\ _06821_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[194]$_DFFE_PP0N_  clock_i _00265_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[14]\ _06820_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[195]$_DFFE_PP0N_  clock_i _00266_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[15]\ _06819_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[196]$_DFFE_PP0N_  clock_i _00267_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[16]\ _06818_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[197]$_DFFE_PP0N_  clock_i _00268_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2101_o[17]\ _06817_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[198]$_DFFE_PP0N_  clock_i _00269_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ _06816_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[199]$_DFFE_PP0N_  clock_i _00270_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _06815_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[19]$_DFFE_PP0N_  clock_i _00271_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[20]\ _06814_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[1]$_DFFE_PP0N_  clock_i _00272_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _06813_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[200]$_DFFE_PP0N_  clock_i _00273_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ _06812_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[201]$_DFFE_PP0N_  clock_i _00274_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _06811_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[202]$_DFFE_PP0N_  clock_i _00275_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ _06810_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[203]$_DFFE_PP0N_  clock_i _00276_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ _06809_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[204]$_DFFE_PP0N_  clock_i _00277_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[6]\ _06808_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[205]$_DFFE_PP0N_  clock_i _00278_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[7]\ _06807_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[206]$_DFFE_PP0N_  clock_i _00279_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[8]\ _06806_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[207]$_DFFE_PP0N_  clock_i _00280_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[9]\ _06805_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[208]$_DFFE_PP0N_  clock_i _00281_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[10]\ _06804_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[209]$_DFFE_PP0N_  clock_i _00282_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[11]\ _06803_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[20]$_DFFE_PP0N_  clock_i _00283_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ _06802_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[210]$_DFFE_PP0N_  clock_i _00284_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[12]\ _06801_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[211]$_DFFE_PP0N_  clock_i _00285_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[13]\ _06800_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[212]$_DFFE_PP0N_  clock_i _00286_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[14]\ _06799_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[213]$_DFFE_PP0N_  clock_i _00287_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[15]\ _06798_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[214]$_DFFE_PP0N_  clock_i _00288_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[16]\ _06797_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[215]$_DFFE_PP0N_  clock_i _00289_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2104_o[17]\ _06796_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[216]$_DFFE_PP0N_  clock_i _00290_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ _06795_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[217]$_DFFE_PP0N_  clock_i _00291_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[229]\ _06794_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[218]$_DFFE_PP0N_  clock_i _00292_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ _06793_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[219]$_DFFE_PP0N_  clock_i _00293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ _06792_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[21]$_DFFE_PP0N_  clock_i _00294_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[22]\ _06791_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[220]$_DFFE_PP0N_  clock_i _00295_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ _06790_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[221]$_DFFE_PP0N_  clock_i _00296_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[233]\ _06789_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[222]$_DFFE_PP0N_  clock_i _00297_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[6]\ _06788_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[223]$_DFFE_PP0N_  clock_i _00298_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[7]\ _06787_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[224]$_DFFE_PP0N_  clock_i _00299_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[8]\ _06786_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[225]$_DFFE_PP0N_  clock_i _00300_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[9]\ _06785_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[226]$_DFFE_PP0N_  clock_i _00301_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[10]\ _06784_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[227]$_DFFE_PP0N_  clock_i _00302_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[11]\ _06783_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[228]$_DFFE_PP0N_  clock_i _00303_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[12]\ _06782_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[229]$_DFFE_PP0N_  clock_i _00304_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[13]\ _06781_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[22]$_DFFE_PP0N_  clock_i _00305_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ _06780_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[230]$_DFFE_PP0N_  clock_i _00306_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[14]\ _06779_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[231]$_DFFE_PP0N_  clock_i _00307_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[15]\ _06778_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[232]$_DFFE_PP0N_  clock_i _00308_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[16]\ _06777_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[233]$_DFFE_PP0N_  clock_i _00309_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2107_o[17]\ _06776_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[234]$_DFFE_PP0N_  clock_i _00310_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ _06775_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[235]$_DFFE_PP0N_  clock_i _00311_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[248]\ _06774_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[236]$_DFFE_PP0N_  clock_i _00312_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ _06773_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[237]$_DFFE_PP0N_  clock_i _00313_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ _06772_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[238]$_DFFE_PP0N_  clock_i _00314_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ _06771_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[239]$_DFFE_PP0N_  clock_i _00315_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[252]\ _06770_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[23]$_DFFE_PP0N_  clock_i _00316_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[24]\ _06769_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[240]$_DFFE_PP0N_  clock_i _00317_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[6]\ _06768_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[241]$_DFFE_PP0N_  clock_i _00318_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[7]\ _06767_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[242]$_DFFE_PP0N_  clock_i _00319_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[8]\ _06766_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[243]$_DFFE_PP0N_  clock_i _00320_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[9]\ _06765_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[244]$_DFFE_PP0N_  clock_i _00321_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[10]\ _06764_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[245]$_DFFE_PP0N_  clock_i _00322_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[11]\ _06763_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[246]$_DFFE_PP0N_  clock_i _00323_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[12]\ _06762_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[247]$_DFFE_PP0N_  clock_i _00324_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[13]\ _06761_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[248]$_DFFE_PP0N_  clock_i _00325_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[14]\ _06760_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[249]$_DFFE_PP0N_  clock_i _00326_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[15]\ _06759_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[24]$_DFFE_PP0N_  clock_i _00327_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[6]\ _06758_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[250]$_DFFE_PP0N_  clock_i _00328_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[16]\ _06757_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[251]$_DFFE_PP0N_  clock_i _00329_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2110_o[17]\ _06756_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[252]$_DFFE_PP0N_  clock_i _00330_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ _06755_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[253]$_DFFE_PP0N_  clock_i _00331_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ _06754_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[254]$_DFFE_PP0N_  clock_i _00332_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ _06753_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[255]$_DFFE_PP0N_  clock_i _00333_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ _06752_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[256]$_DFFE_PP0N_  clock_i _00334_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _06751_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[257]$_DFFE_PP0N_  clock_i _00335_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _06750_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[258]$_DFFE_PP0N_  clock_i _00336_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[6]\ _06749_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[259]$_DFFE_PP0N_  clock_i _00337_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[7]\ _06748_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[25]$_DFFE_PP0N_  clock_i _00338_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[7]\ _06747_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[260]$_DFFE_PP0N_  clock_i _00339_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[8]\ _06746_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[261]$_DFFE_PP0N_  clock_i _00340_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[9]\ _06745_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[262]$_DFFE_PP0N_  clock_i _00341_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[10]\ _06744_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[263]$_DFFE_PP0N_  clock_i _00342_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[11]\ _06743_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[264]$_DFFE_PP0N_  clock_i _00343_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[12]\ _06742_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[265]$_DFFE_PP0N_  clock_i _00344_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[13]\ _06741_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[266]$_DFFE_PP0N_  clock_i _00345_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[14]\ _06740_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[267]$_DFFE_PP0N_  clock_i _00346_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[15]\ _06739_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[268]$_DFFE_PP0N_  clock_i _00347_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[16]\ _06738_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[269]$_DFFE_PP0N_  clock_i _00348_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2443_o[17]\ _06737_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[26]$_DFFE_PP0N_  clock_i _00349_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[8]\ _06736_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[27]$_DFFE_PP0N_  clock_i _00350_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[9]\ _06735_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[28]$_DFFE_PP0N_  clock_i _00351_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[10]\ _06734_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[29]$_DFFE_PP0N_  clock_i _00352_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[11]\ _06733_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[2]$_DFFE_PP0N_  clock_i _00353_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[2]\ _06732_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[30]$_DFFE_PP0N_  clock_i _00354_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[12]\ _06731_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[31]$_DFFE_PP0N_  clock_i _00355_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[13]\ _06730_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[32]$_DFFE_PP0N_  clock_i _00356_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[14]\ _06729_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[33]$_DFFE_PP0N_  clock_i _00357_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[15]\ _06728_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[34]$_DFFE_PP0N_  clock_i _00358_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[16]\ _06727_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[35]$_DFFE_PP0N_  clock_i _00359_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2074_o[17]\ _06726_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[36]$_DFFE_PP0N_  clock_i _00360_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ _06725_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[37]$_DFFE_PP0N_  clock_i _00361_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _06724_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[38]$_DFFE_PP0N_  clock_i _00362_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[40]\ _06723_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[39]$_DFFE_PP0N_  clock_i _00363_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _06722_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[3]$_DFFE_PP0N_  clock_i _00364_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _06721_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[40]$_DFFE_PP0N_  clock_i _00365_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[42]\ _06720_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[41]$_DFFE_PP0N_  clock_i _00366_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[43]\ _06719_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[42]$_DFFE_PP0N_  clock_i _00367_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[6]\ _06718_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[43]$_DFFE_PP0N_  clock_i _00368_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[7]\ _06717_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[44]$_DFFE_PP0N_  clock_i _00369_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[8]\ _06716_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[45]$_DFFE_PP0N_  clock_i _00370_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[9]\ _06715_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[46]$_DFFE_PP0N_  clock_i _00371_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[10]\ _06714_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[47]$_DFFE_PP0N_  clock_i _00372_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[11]\ _06713_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[48]$_DFFE_PP0N_  clock_i _00373_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[12]\ _06712_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[49]$_DFFE_PP0N_  clock_i _00374_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[13]\ _06711_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[4]$_DFFE_PP0N_  clock_i _00375_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[4]\ _06710_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[50]$_DFFE_PP0N_  clock_i _00376_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[14]\ _06709_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[51]$_DFFE_PP0N_  clock_i _00377_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[15]\ _06708_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[52]$_DFFE_PP0N_  clock_i _00378_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[16]\ _06707_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[53]$_DFFE_PP0N_  clock_i _00379_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2077_o[17]\ _06706_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[54]$_DFFE_PP0N_  clock_i _00380_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ _06705_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[55]$_DFFE_PP0N_  clock_i _00381_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[58]\ _06704_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[56]$_DFFE_PP0N_  clock_i _00382_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[59]\ _06703_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[57]$_DFFE_PP0N_  clock_i _00383_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[60]\ _06702_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[58]$_DFFE_PP0N_  clock_i _00384_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ _06701_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[59]$_DFFE_PP0N_  clock_i _00385_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[62]\ _06700_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[5]$_DFFE_PP0N_  clock_i _00386_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ _06699_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[60]$_DFFE_PP0N_  clock_i _00387_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[6]\ _06698_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[61]$_DFFE_PP0N_  clock_i _00388_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[7]\ _06697_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[62]$_DFFE_PP0N_  clock_i _00389_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[8]\ _06696_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[63]$_DFFE_PP0N_  clock_i _00390_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[9]\ _06695_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[64]$_DFFE_PP0N_  clock_i _00391_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[10]\ _06694_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[65]$_DFFE_PP0N_  clock_i _00392_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[11]\ _06693_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[66]$_DFFE_PP0N_  clock_i _00393_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[12]\ _06692_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[67]$_DFFE_PP0N_  clock_i _00394_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[13]\ _06691_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[68]$_DFFE_PP0N_  clock_i _00395_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[14]\ _06690_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[69]$_DFFE_PP0N_  clock_i _00396_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[15]\ _06689_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[6]$_DFFE_PP0N_  clock_i _00397_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[6]\ _06688_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[70]$_DFFE_PP0N_  clock_i _00398_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[16]\ _06687_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[71]$_DFFE_PP0N_  clock_i _00399_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2080_o[17]\ _06686_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[72]$_DFFE_PP0N_  clock_i _00400_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ _06685_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[73]$_DFFE_PP0N_  clock_i _00401_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _06684_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[74]$_DFFE_PP0N_  clock_i _00402_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ _06683_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[75]$_DFFE_PP0N_  clock_i _00403_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _06682_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[76]$_DFFE_PP0N_  clock_i _00404_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _06681_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[77]$_DFFE_PP0N_  clock_i _00405_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[81]\ _06680_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[78]$_DFFE_PP0N_  clock_i _00406_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[6]\ _06679_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[79]$_DFFE_PP0N_  clock_i _00407_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[7]\ _06678_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[7]$_DFFE_PP0N_  clock_i _00408_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[7]\ _06677_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[80]$_DFFE_PP0N_  clock_i _00409_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[8]\ _06676_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[81]$_DFFE_PP0N_  clock_i _00410_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[9]\ _06675_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[82]$_DFFE_PP0N_  clock_i _00411_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[10]\ _06674_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[83]$_DFFE_PP0N_  clock_i _00412_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[11]\ _06673_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[84]$_DFFE_PP0N_  clock_i _00413_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[12]\ _06672_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[85]$_DFFE_PP0N_  clock_i _00414_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[13]\ _06671_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[86]$_DFFE_PP0N_  clock_i _00415_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[14]\ _06670_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[87]$_DFFE_PP0N_  clock_i _00416_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[15]\ _06669_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[88]$_DFFE_PP0N_  clock_i _00417_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[16]\ _06668_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[89]$_DFFE_PP0N_  clock_i _00418_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2083_o[17]\ _06667_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[8]$_DFFE_PP0N_  clock_i _00419_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[8]\ _06666_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[90]$_DFFE_PP0N_  clock_i _00420_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ _06665_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[91]$_DFFE_PP0N_  clock_i _00421_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ _06664_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[92]$_DFFE_PP0N_  clock_i _00422_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ _06663_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[93]$_DFFE_PP0N_  clock_i _00423_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ _06662_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[94]$_DFFE_PP0N_  clock_i _00424_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ _06661_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[95]$_DFFE_PP0N_  clock_i _00425_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _06660_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[96]$_DFFE_PP0N_  clock_i _00426_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[6]\ _06659_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[97]$_DFFE_PP0N_  clock_i _00427_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[7]\ _06658_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[98]$_DFFE_PP0N_  clock_i _00428_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[8]\ _06657_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[99]$_DFFE_PP0N_  clock_i _00429_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2086_o[9]\ _06656_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2459_q[9]$_DFFE_PP0N_  clock_i _00430_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2071_o[9]\ _06655_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[0]$_DFFE_PP0P_  clock_i _00431_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2070_o[0]\ _00089_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[10]$_DFFE_PP0P_  clock_i _00432_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2085_o[0]\ _00080_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[11]$_DFFE_PP0P_  clock_i _00433_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2085_o[1]\ _06654_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[12]$_DFFE_PP0P_  clock_i _00434_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2088_o[0]\ _06653_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[13]$_DFFE_PP0P_  clock_i _00435_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2088_o[1]\ _06652_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[14]$_DFFE_PP0P_  clock_i _00436_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2091_o[0]\ _06651_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[15]$_DFFE_PP0P_  clock_i _00437_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2091_o[1]\ _06650_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[16]$_DFFE_PP0P_  clock_i _00438_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2094_o[0]\ _00076_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[17]$_DFFE_PP0P_  clock_i _00439_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2094_o[1]\ _06649_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[18]$_DFFE_PP0P_  clock_i _00440_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2097_o[0]\ _00075_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[19]$_DFFE_PP0P_  clock_i _00441_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2097_o[1]\ _06648_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[1]$_DFFE_PP0P_  clock_i _00442_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2070_o[1]\ _06647_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[20]$_DFFE_PP0P_  clock_i _00443_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2100_o[0]\ _00074_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[21]$_DFFE_PP0P_  clock_i _00444_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2100_o[1]\ _06646_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[22]$_DFFE_PP0P_  clock_i _00445_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2103_o[0]\ _00071_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[23]$_DFFE_PP0P_  clock_i _00446_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2103_o[1]\ _06645_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[24]$_DFFE_PP0P_  clock_i _00447_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2106_o[0]\ _00072_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[25]$_DFFE_PP0P_  clock_i _00448_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2106_o[1]\ _06644_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[26]$_DFFE_PP0P_  clock_i _00449_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2109_o[0]\ _00073_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[27]$_DFFE_PP0P_  clock_i _00450_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2109_o[1]\ _06643_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[28]$_DFFE_PP0P_  clock_i _00451_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2934_o\ _06642_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[29]$_DFFE_PP0P_  clock_i _00452_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n2931_o\ _06641_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[2]$_DFFE_PP0P_  clock_i _00453_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2073_o[0]\ _00088_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[3]$_DFFE_PP0P_  clock_i _00454_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2073_o[1]\ _06640_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[4]$_DFFE_PP0P_  clock_i _00455_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2076_o[0]\ _00086_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[5]$_DFFE_PP0P_  clock_i _00456_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2076_o[1]\ _06639_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[6]$_DFFE_PP0P_  clock_i _00457_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2079_o[0]\ _00084_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[7]$_DFFE_PP0P_  clock_i _00458_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2079_o[1]\ _06638_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[8]$_DFFE_PP0P_  clock_i _00459_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2082_o[0]\ _00082_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2460_q[9]$_DFFE_PP0P_  clock_i _00460_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2082_o[1]\ _06637_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[0]$_DFFE_PP0P_  clock_i _00461_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2072_o\ _06636_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[10]$_DFFE_PP0P_  clock_i _00462_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2102_o\ _06635_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[11]$_DFFE_PP0P_  clock_i _00463_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2105_o\ _06634_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[12]$_DFFE_PP0P_  clock_i _00464_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2108_o\ _06633_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[13]$_DFFE_PP0P_  clock_i _00465_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2111_o\ _06632_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[14]$_DFFE_PP0P_  clock_i _00466_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2446_o\ _06631_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[1]$_DFFE_PP0P_  clock_i _00467_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2075_o\ _06630_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[2]$_DFFE_PP0P_  clock_i _00468_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2078_o\ _06629_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[3]$_DFFE_PP0P_  clock_i _00469_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2081_o\ _06628_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[4]$_DFFE_PP0P_  clock_i _00470_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2084_o\ _06627_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[5]$_DFFE_PP0P_  clock_i _00471_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2087_o\ _06626_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[6]$_DFFE_PP0P_  clock_i _00472_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2090_o\ _06625_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[7]$_DFFE_PP0P_  clock_i _00473_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2093_o\ _06624_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[8]$_DFFE_PP0P_  clock_i _00474_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2096_o\ _06623_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2462_q[9]$_DFFE_PP0P_  clock_i _00475_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2099_o\ _06622_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2463_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2213_o\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2463_q\ _06621_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[48]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[0]\ _00079_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[49]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ _00081_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[2]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[50]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ _00083_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[3]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[51]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _00085_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[4]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[52]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ _00087_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2671_q[5]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[53]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _06620_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2672_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1321_o\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2468_o\ _06619_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2672_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2468_o\ \atbs_core_0.adaptive_ctrl_0.n1352_o\ _00051_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[0]\ _06618_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[1]\ _06617_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[2]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2669_o[2]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n2677_q[2]\ _06616_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1585_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1498_o\ \atbs_core_0.dac_control_0.n1495_o\ _00028_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1586_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1495_o\ \atbs_core_0.dac_control_0.n1586_q\ _00047_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[1]$_DFFE_PP0N_  clock_i _00476_ \atbs_core_0.dac_control_0.dac_init_value[1]\ _06615_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[2]$_DFFE_PP0N_  clock_i _00477_ \atbs_core_0.dac_control_0.dac_init_value[2]\ _06614_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[3]$_DFFE_PP0N_  clock_i _00478_ \atbs_core_0.dac_control_0.dac_init_value[3]\ _06613_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[4]$_DFFE_PP0N_  clock_i _00479_ \atbs_core_0.dac_control_0.dac_init_value[4]\ _06612_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[5]$_DFFE_PP0N_  clock_i _00480_ \atbs_core_0.dac_control_0.dac_init_value[5]\ _06611_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[6]$_DFFE_PP0N_  clock_i _00481_ \atbs_core_0.dac_control_0.dac_init_value[6]\ _06610_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[7]$_DFFE_PP0N_  clock_i _00482_ \atbs_core_0.dac_control_0.dac_init_value[7]\ _06609_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1587_q[8]$_DFFE_PP0N_  clock_i _00483_ \atbs_core_0.dac_control_0.dac_init_value[8]\ _06608_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[0]$_DFFE_PP0P_  clock_i _00484_ \atbs_core_0.dac_control_0.dac_counter_value[0]\ _00069_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[1]$_DFFE_PP0P_  clock_i _00485_ \atbs_core_0.dac_control_0.dac_counter_value[1]\ _00044_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[2]$_DFFE_PP0P_  clock_i _00486_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ _00042_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[3]$_DFFE_PP0P_  clock_i _00487_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ _00041_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[4]$_DFFE_PP0P_  clock_i _00488_ \atbs_core_0.dac_control_0.dac_counter_value[4]\ _00038_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[5]$_DFFE_PP0P_  clock_i _00489_ \atbs_core_0.dac_control_0.dac_counter_value[5]\ _00037_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[6]$_DFFE_PP0P_  clock_i _00490_ \atbs_core_0.dac_control_0.dac_counter_value[6]\ _06607_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[7]$_DFFE_PP0P_  clock_i _00491_ \atbs_core_0.dac_control_0.dac_counter_value[7]\ _06606_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1588_q[8]$_DFFE_PP0P_  clock_i _00492_ \atbs_core_0.dac_control_0.dac_counter_value[8]\ _00070_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[0]$_DFFE_PP0P_  clock_i _00493_ dac_upper_o[0] _06605_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[1]$_DFFE_PP0P_  clock_i _00494_ dac_upper_o[1] _06604_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[2]$_DFFE_PP0P_  clock_i _00495_ dac_upper_o[2] _06603_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[3]$_DFFE_PP0P_  clock_i _00496_ dac_upper_o[3] _06602_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[4]$_DFFE_PP0P_  clock_i _00497_ dac_upper_o[4] _00078_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[5]$_DFFE_PP0P_  clock_i _00498_ dac_upper_o[5] _06601_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[6]$_DFFE_PP0P_  clock_i _00499_ dac_upper_o[6] _06600_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1590_q[7]$_DFFE_PP0P_  clock_i _00500_ dac_upper_o[7] _06599_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1591_q$_DFFE_PP0P_  clock_i _00501_ \atbs_core_0.dac_control_0.dac_change_in_progress\ _06598_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1592_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1566_o[0]\ \atbs_core_0.dac_control_0.n1592_q[0]\ _06597_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1592_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1566_o[1]\ \atbs_core_0.dac_control_0.n1592_q[1]\ _06596_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1592_q[2]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1566_o[2]\ \atbs_core_0.dac_control_0.n1592_q[2]\ _00030_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.dac_counter_strb\ \atbs_core_0.dac_control_0.sync_chain_0.n1088_o\ _06595_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.sync_chain_0.n1088_o\ \atbs_core_0.dac_control_0.dac_wr_o\ _06594_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1720_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1632_o\ \atbs_core_0.dac_control_1.n1629_o\ _06593_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1721_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1629_o\ \atbs_core_0.dac_control_1.n1721_q\ _00054_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1722_q[7]$_DFFE_PP0N_  clock_i _00502_ \atbs_core_0.dac_control_1.dac_init_value[7]\ _06592_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[0]$_DFFE_PP0P_  clock_i _00503_ \atbs_core_0.dac_control_1.dac_counter_value[0]\ _00067_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[1]$_DFFE_PP0P_  clock_i _00504_ \atbs_core_0.dac_control_1.dac_counter_value[1]\ _00059_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[2]$_DFFE_PP0P_  clock_i _00505_ \atbs_core_0.dac_control_1.dac_counter_value[2]\ _00058_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[3]$_DFFE_PP0P_  clock_i _00506_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ _00057_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[4]$_DFFE_PP0P_  clock_i _00507_ \atbs_core_0.dac_control_1.dac_counter_value[4]\ _00056_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[5]$_DFFE_PP0P_  clock_i _00508_ \atbs_core_0.dac_control_1.dac_counter_value[5]\ _00055_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[6]$_DFFE_PP0P_  clock_i _00509_ \atbs_core_0.dac_control_1.dac_counter_value[6]\ _06591_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[7]$_DFFE_PP0P_  clock_i _00510_ \atbs_core_0.dac_control_1.dac_counter_value[7]\ _06590_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1723_q[8]$_DFFE_PP0P_  clock_i _00511_ \atbs_core_0.dac_control_1.dac_counter_value[8]\ _00068_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[0]$_DFFE_PP0P_  clock_i _00512_ dac_lower_o[0] _06589_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[1]$_DFFE_PP0P_  clock_i _00513_ dac_lower_o[1] _06588_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[2]$_DFFE_PP0P_  clock_i _00514_ dac_lower_o[2] _06587_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[3]$_DFFE_PP0P_  clock_i _00515_ dac_lower_o[3] _06586_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[4]$_DFFE_PP0P_  clock_i _00516_ dac_lower_o[4] _06585_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[5]$_DFFE_PP0P_  clock_i _00517_ dac_lower_o[5] _06584_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[6]$_DFFE_PP0P_  clock_i _00518_ dac_lower_o[6] _06583_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1725_q[7]$_DFFE_PP0P_  clock_i _00519_ dac_lower_o[7] _06582_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1726_q$_DFFE_PP0P_  clock_i _00520_ \atbs_core_0.dac_control_1.dac_change_in_progress\ _06581_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1727_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1701_o[0]\ \atbs_core_0.dac_control_1.n1727_q[0]\ _06580_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1727_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1701_o[1]\ \atbs_core_0.dac_control_1.n1727_q[1]\ _06579_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n1727_q[2]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1701_o[2]\ \atbs_core_0.dac_control_1.n1727_q[2]\ _00053_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.dac_counter_strb\ \atbs_core_0.dac_control_1.sync_chain_0.n1088_o\ _06578_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.sync_chain_0.n1088_o\ \atbs_core_0.dac_control_1.dac_wr_o\ _06577_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.bouncing_sync\ \atbs_core_0.debouncer_0.bouncing_sync_d\ _06576_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1128_o[0]\ \atbs_core_0.debouncer_0.counter_value[0]\ _06575_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1128_o[1]\ \atbs_core_0.debouncer_0.counter_value[1]\ _06574_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1128_o[2]\ \atbs_core_0.debouncer_0.counter_value[2]\ _06573_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1128_o[3]\ \atbs_core_0.debouncer_0.counter_value[3]\ _06572_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1173_q[0]$_DFFE_PP0P_  clock_i _00521_ \atbs_core_0.debouncer_0.n1173_q[0]\ _06571_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1173_q[1]$_DFFE_PP0P_  clock_i _00522_ \atbs_core_0.debouncer_0.n1173_q[1]\ _06570_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1174_q$_DFFE_PP0P_  clock_i _00523_ \atbs_core_0.debouncer_0.debounced\ _06569_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i trigger_start_mode_i \atbs_core_0.debouncer_0.sync_chain_0.n1088_o\ _06568_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_0.bouncing_sync\ _06567_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.bouncing_sync\ \atbs_core_0.debouncer_1.bouncing_sync_d\ _06566_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1128_o[0]\ \atbs_core_0.debouncer_1.counter_value[0]\ _06565_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1128_o[1]\ \atbs_core_0.debouncer_1.counter_value[1]\ _06564_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1128_o[2]\ \atbs_core_0.debouncer_1.counter_value[2]\ _06563_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1128_o[3]\ \atbs_core_0.debouncer_1.counter_value[3]\ _06562_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1173_q[0]$_DFFE_PP0P_  clock_i _00524_ \atbs_core_0.debouncer_1.n1173_q[0]\ _06561_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1173_q[1]$_DFFE_PP0P_  clock_i _00525_ \atbs_core_0.debouncer_1.n1173_q[1]\ _06560_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1174_q$_DFFE_PP0P_  clock_i _00526_ \atbs_core_0.adaptive_mode_debounced\ _00008_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i adaptive_mode_i \atbs_core_0.debouncer_1.sync_chain_0.n1088_o\ _06559_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_1.bouncing_sync\ _06558_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.bouncing_sync\ \atbs_core_0.debouncer_2.bouncing_sync_d\ _06557_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1128_o[0]\ \atbs_core_0.debouncer_2.counter_value[0]\ _06556_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1128_o[1]\ \atbs_core_0.debouncer_2.counter_value[1]\ _06555_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1128_o[2]\ \atbs_core_0.debouncer_2.counter_value[2]\ _06554_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1128_o[3]\ \atbs_core_0.debouncer_2.counter_value[3]\ _06553_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1173_q[0]$_DFFE_PP0P_  clock_i _00527_ \atbs_core_0.debouncer_2.n1173_q[0]\ _06552_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1173_q[1]$_DFFE_PP0P_  clock_i _00528_ \atbs_core_0.debouncer_2.n1173_q[1]\ _06551_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1174_q$_DFFE_PP0P_  clock_i _00529_ \atbs_core_0.control_mode_debounced\ _06550_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i control_mode_i \atbs_core_0.debouncer_2.sync_chain_0.n1088_o\ _06549_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_2.bouncing_sync\ _06548_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.bouncing_sync\ \atbs_core_0.debouncer_3.bouncing_sync_d\ _06547_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1128_o[0]\ \atbs_core_0.debouncer_3.counter_value[0]\ _06546_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1128_o[1]\ \atbs_core_0.debouncer_3.counter_value[1]\ _06545_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1128_o[2]\ \atbs_core_0.debouncer_3.counter_value[2]\ _06544_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1128_o[3]\ \atbs_core_0.debouncer_3.counter_value[3]\ _06543_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1173_q[0]$_DFFE_PP0P_  clock_i _00530_ \atbs_core_0.debouncer_3.n1173_q[0]\ _06542_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1173_q[1]$_DFFE_PP0P_  clock_i _00531_ \atbs_core_0.debouncer_3.n1173_q[1]\ _06541_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1174_q$_DFFE_PP0P_  clock_i _00532_ \atbs_core_0.debouncer_3.debounced\ _06540_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i signal_select_in_i \atbs_core_0.debouncer_3.sync_chain_0.n1088_o\ _06539_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_3.bouncing_sync\ _06538_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.bouncing_sync\ \atbs_core_0.debouncer_4.bouncing_sync_d\ _06537_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1128_o[0]\ \atbs_core_0.debouncer_4.counter_value[0]\ _06536_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1128_o[1]\ \atbs_core_0.debouncer_4.counter_value[1]\ _06535_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1128_o[2]\ \atbs_core_0.debouncer_4.counter_value[2]\ _06534_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1128_o[3]\ \atbs_core_0.debouncer_4.counter_value[3]\ _06533_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1173_q[0]$_DFFE_PP0P_  clock_i _00533_ \atbs_core_0.debouncer_4.n1173_q[0]\ _06532_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1173_q[1]$_DFFE_PP0P_  clock_i _00534_ \atbs_core_0.debouncer_4.n1173_q[1]\ _06531_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1174_q$_DFFE_PP0P_  clock_i _00535_ \atbs_core_0.debouncer_4.debounced\ _06530_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i enable_i \atbs_core_0.debouncer_4.sync_chain_0.n1088_o\ _06529_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_4.bouncing_sync\ _06528_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1171_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.bouncing_sync\ \atbs_core_0.debouncer_5.bouncing_sync_d\ _06527_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1172_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1128_o[0]\ \atbs_core_0.debouncer_5.counter_value[0]\ _06526_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1172_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1128_o[1]\ \atbs_core_0.debouncer_5.counter_value[1]\ _06525_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1172_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1128_o[2]\ \atbs_core_0.debouncer_5.counter_value[2]\ _06524_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1172_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1128_o[3]\ \atbs_core_0.debouncer_5.counter_value[3]\ _06523_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1173_q[0]$_DFFE_PP0P_  clock_i _00536_ \atbs_core_0.debouncer_5.n1173_q[0]\ _06522_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1173_q[1]$_DFFE_PP0P_  clock_i _00537_ \atbs_core_0.debouncer_5.n1173_q[1]\ _06521_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1174_q$_DFFE_PP0P_  clock_i _00538_ \atbs_core_0.debouncer_5.debounced\ _06520_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.sync_chain_0.n1095_q[0]$_DFF_PP0_  clock_i select_tbs_delta_steps_i \atbs_core_0.debouncer_5.sync_chain_0.n1088_o\ _06519_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.sync_chain_0.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.sync_chain_0.n1088_o\ \atbs_core_0.debouncer_5.bouncing_sync\ _06518_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[0]$_DFFE_PP0P_  clock_i _00539_ \atbs_core_0.uart_0.uart_tx_0.n2783_o\ _06517_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[10]$_DFFE_PP0P_  clock_i _00540_ \atbs_core_0.memory2uart_0.n2009_o[2]\ _06516_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[11]$_DFFE_PP0P_  clock_i _00541_ \atbs_core_0.memory2uart_0.n2009_o[3]\ _06515_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[12]$_DFFE_PP0P_  clock_i _00542_ \atbs_core_0.memory2uart_0.n2009_o[4]\ _06514_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[13]$_DFFE_PP0P_  clock_i _00543_ \atbs_core_0.memory2uart_0.n2009_o[5]\ _06513_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[14]$_DFFE_PP0P_  clock_i _00544_ \atbs_core_0.memory2uart_0.n2009_o[6]\ _06512_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[15]$_DFFE_PP0P_  clock_i _00545_ \atbs_core_0.memory2uart_0.n2009_o[7]\ _06511_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[16]$_DFFE_PP0P_  clock_i _00546_ \atbs_core_0.memory2uart_0.n2009_o[8]\ _06510_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[17]$_DFFE_PP0P_  clock_i _00547_ \atbs_core_0.memory2uart_0.n2009_o[9]\ _06509_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[18]$_DFFE_PP0P_  clock_i _00548_ \atbs_core_0.memory2uart_0.n2009_o[10]\ _06508_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[19]$_DFFE_PP0P_  clock_i _00549_ \atbs_core_0.memory2uart_0.n2009_o[11]\ _06507_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[1]$_DFFE_PP0P_  clock_i _00550_ \atbs_core_0.uart_0.uart_tx_0.n2784_o\ _06506_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[20]$_DFFE_PP0P_  clock_i _00551_ \atbs_core_0.memory2uart_0.n2009_o[12]\ _06505_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[21]$_DFFE_PP0P_  clock_i _00552_ \atbs_core_0.memory2uart_0.n2009_o[13]\ _06504_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[22]$_DFFE_PP0P_  clock_i _00553_ \atbs_core_0.memory2uart_0.n2009_o[14]\ _06503_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[23]$_DFFE_PP0P_  clock_i _00554_ \atbs_core_0.memory2uart_0.n2009_o[15]\ _06502_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[2]$_DFFE_PP0P_  clock_i _00555_ \atbs_core_0.uart_0.uart_tx_0.n2785_o\ _06501_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[3]$_DFFE_PP0P_  clock_i _00556_ \atbs_core_0.uart_0.uart_tx_0.n2786_o\ _06500_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[4]$_DFFE_PP0P_  clock_i _00557_ \atbs_core_0.uart_0.uart_tx_0.n2787_o\ _06499_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[5]$_DFFE_PP0P_  clock_i _00558_ \atbs_core_0.uart_0.uart_tx_0.n2788_o\ _06498_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[6]$_DFFE_PP0P_  clock_i _00559_ \atbs_core_0.uart_0.uart_tx_0.n2789_o\ _06497_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[7]$_DFFE_PP0P_  clock_i _00560_ \atbs_core_0.uart_0.uart_tx_0.n2790_o\ _06496_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[8]$_DFFE_PP0P_  clock_i _00561_ \atbs_core_0.memory2uart_0.n2009_o[0]\ _06495_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2038_q[9]$_DFFE_PP0P_  clock_i _00562_ \atbs_core_0.memory2uart_0.n2009_o[1]\ _06494_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2040_q$_DFF_PP0_  clock_i \atbs_core_0.memory2uart_0.n2023_o\ \atbs_core_0.memory2uart_0.n2040_q\ _00031_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2041_q[0]$_DFFE_PP0P_  clock_i _00563_ \atbs_core_0.memory2uart_0.counter[0]\ _06493_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2041_q[1]$_DFFE_PP0P_  clock_i _00564_ \atbs_core_0.memory2uart_0.counter[1]\ _06492_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1046_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_mode_debounced\ \atbs_core_0.adaptive_mode_d\ _06491_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1047_q$_DFF_PP0_  clock_i \atbs_core_0.control_mode_debounced\ \atbs_core_0.control_mode_d\ _06490_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1048_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.debounced\ \atbs_core_0.n1048_q\ _06489_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1049_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.debounced\ \atbs_core_0.n1049_q\ _06488_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1050_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.debounced\ \atbs_core_0.n1050_q\ _06487_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1051_q$_DFF_PP0_  clock_i \atbs_core_0.n37_o\ \atbs_core_0.n1051_q\ _06486_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1052_q$_DFFE_PP0P_  clock_i _00565_ \atbs_core_0.detection_en\ _06485_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1053_q$_DFF_PP0_  clock_i \atbs_core_0.n148_o\ \atbs_core_0.n1053_q\ _06484_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1054_q$_DFF_PP0_  clock_i \atbs_core_0.n156_o\ \atbs_core_0.n1054_q\ _06483_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1056_q$_DFFE_PP0P_  clock_i _00566_ \atbs_core_0.n1056_q\ _06482_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1057_q$_DFFE_PP0P_  clock_i _00567_ \atbs_core_0.enable_read\ _06481_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1058_q$_DFFE_PP0P_  clock_i _00568_ \atbs_core_0.analog_trigger_uart\ _00050_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1061_q$_DFFE_PP0P_  clock_i _00569_ \atbs_core_0.n1061_q\ _06480_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1065_q$_DFFE_PP0P_  clock_i _00570_ \atbs_core_0.baudrate_uart\ _00048_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[0]$_DFFE_PP1P_  clock_i _00571_ _00105_ \atbs_core_0.baudrate_adj_uart[0]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[2]$_DFFE_PP1P_  clock_i _00572_ _00106_ \atbs_core_0.baudrate_adj_uart[2]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[3]$_DFFE_PP0P_  clock_i _00573_ \atbs_core_0.baudrate_adj_uart[1]\ _06479_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[4]$_DFFE_PP0P_  clock_i _00574_ \atbs_core_0.baudrate_adj_uart[4]\ _06478_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[5]$_DFFE_PP0P_  clock_i _00575_ \atbs_core_0.baudrate_adj_uart[5]\ _06477_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[6]$_DFFE_PP1P_  clock_i _00576_ _00107_ \atbs_core_0.baudrate_adj_uart[6]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1066_q[7]$_DFFE_PP0P_  clock_i _00577_ \atbs_core_0.baudrate_adj_uart[7]\ _06476_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1067_q$_DFFE_PP0P_  clock_i _00578_ \atbs_core_0.n1067_q\ _00049_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1068_q[1]$_DFFE_PP0P_  clock_i _00579_ \atbs_core_0.n1068_q[1]\ _06475_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1068_q[2]$_DFFE_PP0P_  clock_i _00580_ \atbs_core_0.n1068_q[2]\ _06474_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1068_q[3]$_DFFE_PP1P_  clock_i _00581_ _00108_ \atbs_core_0.n1068_q[3]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1068_q[4]$_DFFE_PP0P_  clock_i _00582_ \atbs_core_0.n1068_q[4]\ _06473_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1068_q[5]$_DFFE_PP0P_  clock_i _00583_ \atbs_core_0.n1068_q[5]\ _06472_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1069_q$_DFFE_PP0P_  clock_i _00584_ \atbs_core_0.atbs_win_length_uart\ _06471_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[10]$_DFFE_PP1P_  clock_i _00585_ _00109_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[10]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[11]$_DFFE_PP1P_  clock_i _00586_ _00110_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[11]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[12]$_DFFE_PP1P_  clock_i _00587_ _00111_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[12]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[13]$_DFFE_PP1P_  clock_i _00588_ _00112_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[13]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[14]$_DFFE_PP1P_  clock_i _00589_ _00113_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[14]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[15]$_DFFE_PP0P_  clock_i _00590_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[15]\ _06470_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[16]$_DFFE_PP0P_  clock_i _00591_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[16]\ _06469_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[17]$_DFFE_PP0P_  clock_i _00592_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[17]\ _06468_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[6]$_DFFE_PP0P_  clock_i _00593_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[6]\ _06467_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[7]$_DFFE_PP0P_  clock_i _00594_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[7]\ _06466_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[8]$_DFFE_PP1P_  clock_i _00595_ _00114_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[8]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1070_q[9]$_DFFE_PP0P_  clock_i _00596_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[9]\ _06465_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1071_q$_DFFE_PP0P_  clock_i _00597_ \atbs_core_0.atbs_max_delta_steps_uart\ _00077_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1072_q[2]$_DFFE_PP0P_  clock_i _00598_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _06464_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1072_q[3]$_DFFE_PP0P_  clock_i _00599_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _06463_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1072_q[4]$_DFFE_PP0P_  clock_i _00600_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _06462_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1072_q[5]$_DFFE_PP1P_  clock_i _00601_ _00115_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[5]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1072_q[6]$_DFFE_PP0P_  clock_i _00602_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[6]\ _06461_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[0]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[0]\ \atbs_core_0.main_counter_value[0]\ _06460_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[10]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[10]\ \atbs_core_0.main_counter_value[10]\ _06459_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[11]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[11]\ \atbs_core_0.main_counter_value[11]\ _06458_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[12]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[12]\ \atbs_core_0.main_counter_value[12]\ _06457_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[13]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[13]\ \atbs_core_0.main_counter_value[13]\ _06456_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[14]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[14]\ \atbs_core_0.main_counter_value[14]\ _06455_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[15]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[15]\ \atbs_core_0.main_counter_value[15]\ _06454_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[16]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[16]\ \atbs_core_0.main_counter_value[16]\ _06453_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[17]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[17]\ \atbs_core_0.main_counter_value[17]\ _06452_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[18]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[18]\ \atbs_core_0.main_counter_value[18]\ _06451_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[19]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[19]\ \atbs_core_0.main_counter_value[19]\ _06450_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[1]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[1]\ \atbs_core_0.main_counter_value[1]\ _06449_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[2]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[2]\ \atbs_core_0.main_counter_value[2]\ _06448_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[3]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[3]\ \atbs_core_0.main_counter_value[3]\ _06447_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[4]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[4]\ \atbs_core_0.main_counter_value[4]\ _06446_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[5]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[5]\ \atbs_core_0.main_counter_value[5]\ _06445_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[6]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[6]\ \atbs_core_0.main_counter_value[6]\ _06444_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[7]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[7]\ \atbs_core_0.main_counter_value[7]\ _06443_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[8]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[8]\ \atbs_core_0.main_counter_value[8]\ _06442_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1073_q[9]$_DFF_PP0_  clock_i \atbs_core_0.n206_o[9]\ \atbs_core_0.main_counter_value[9]\ _06441_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1074_q[0]$_DFF_PP1_  clock_i _00121_ _06937_ \atbs_core_0.n1074_q[0]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1074_q[1]$_DFF_PP0_  clock_i \atbs_core_0.n391_o[1]\ \atbs_core_0.n1074_q[1]\ _06440_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1074_q[2]$_DFF_PP0_  clock_i \atbs_core_0.n391_o[2]\ \atbs_core_0.n1074_q[2]\ _00027_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1075_q$_DFFE_PP0P_  clock_i _00603_ idle_led_o _06439_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1076_q$_DFFE_PP0P_  clock_i _00604_ overflow_led_o _06438_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1077_q$_DFFE_PP0P_  clock_i _00605_ underflow_led_o _06437_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1078_q$_DFFE_PP1P_  clock_i _00606_ _00116_ \atbs_core_0.n1078_q\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1079_q$_DFFE_PP0P_  clock_i _00607_ \atbs_core_0.adaptive_mode_uart\ _00009_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1081_q$_DFFE_PP1P_  clock_i _00608_ _00117_ \atbs_core_0.enable_analog_uart\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1082_q$_DFFE_PP1P_  clock_i _00609_ _00118_ \atbs_core_0.n1082_q\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1256_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.spike_i\ \atbs_core_0.spike_detector_0.hold_spike\ _00025_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1257_q$_DFFE_PP0P_  clock_i _00610_ \atbs_core_0.spike_detector_0.lock_detection\ _06436_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1258_q$_DFFE_PP0P_  clock_i _00611_ \atbs_core_0.spike_detector_0.n1258_q\ _06435_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1259_q$_DFFE_PP0P_  clock_i _00612_ \atbs_core_0.spike_detector_0.lower_is_changing\ _06434_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1260_q$_DFF_PP0_  clock_i \atbs_core_0.spike_detector_0.n1246_o\ \atbs_core_0.spike_detector_0.is_changing\ _06433_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[0]$_DFFE_PP0P_  clock_i _00613_ \atbs_core_0.encoded_spike[0]\ _06432_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[10]$_DFFE_PP0P_  clock_i _00614_ \atbs_core_0.encoded_spike[10]\ _06431_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[11]$_DFFE_PP0P_  clock_i _00615_ \atbs_core_0.encoded_spike[11]\ _06430_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[12]$_DFFE_PP0P_  clock_i _00616_ \atbs_core_0.encoded_spike[12]\ _06429_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[13]$_DFFE_PP0P_  clock_i _00617_ \atbs_core_0.encoded_spike[13]\ _06428_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[14]$_DFFE_PP0P_  clock_i _00618_ \atbs_core_0.encoded_spike[14]\ _06427_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[15]$_DFFE_PP0P_  clock_i _00619_ \atbs_core_0.encoded_spike[15]\ _06426_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[16]$_DFFE_PP0P_  clock_i _00620_ \atbs_core_0.encoded_spike[16]\ _06425_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[17]$_DFFE_PP0P_  clock_i _00621_ \atbs_core_0.encoded_spike[17]\ _06424_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[18]$_DFFE_PP0P_  clock_i _00622_ \atbs_core_0.encoded_spike[18]\ _06423_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[1]$_DFFE_PP0P_  clock_i _00623_ \atbs_core_0.encoded_spike[1]\ _06422_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[2]$_DFFE_PP0P_  clock_i _00624_ \atbs_core_0.encoded_spike[2]\ _06421_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[3]$_DFFE_PP0P_  clock_i _00625_ \atbs_core_0.encoded_spike[3]\ _06420_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[4]$_DFFE_PP0P_  clock_i _00626_ \atbs_core_0.encoded_spike[4]\ _06419_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[5]$_DFFE_PP0P_  clock_i _00627_ \atbs_core_0.encoded_spike[5]\ _06418_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[6]$_DFFE_PP0P_  clock_i _00628_ \atbs_core_0.encoded_spike[6]\ _06417_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[7]$_DFFE_PP0P_  clock_i _00629_ \atbs_core_0.encoded_spike[7]\ _06416_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[8]$_DFFE_PP0P_  clock_i _00630_ \atbs_core_0.encoded_spike[8]\ _06415_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1865_q[9]$_DFFE_PP0P_  clock_i _00631_ \atbs_core_0.encoded_spike[9]\ _06414_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1866_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n1860_o\ \atbs_core_0.encoded_spike_strb\ _06413_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1867_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n1839_o\ \atbs_core_0.spike_encoder_0.delayed_spike_strb\ _06412_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n1868_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n1845_o\ \atbs_core_0.spike_encoder_0.delayed_spike\ _06411_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[0]$_DFFE_PP0P_  clock_i _00632_ \atbs_core_0.spike_memory_0.n1953_o[0]\ _06410_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[10]$_DFFE_PP0P_  clock_i _00633_ \atbs_core_0.spike_memory_0.n1953_o[10]\ _06409_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[11]$_DFFE_PP0P_  clock_i _00634_ \atbs_core_0.spike_memory_0.n1953_o[11]\ _06408_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[12]$_DFFE_PP0P_  clock_i _00635_ \atbs_core_0.spike_memory_0.n1953_o[12]\ _06407_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[13]$_DFFE_PP0P_  clock_i _00636_ \atbs_core_0.spike_memory_0.n1953_o[13]\ _06406_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[14]$_DFFE_PP0P_  clock_i _00637_ \atbs_core_0.spike_memory_0.n1953_o[14]\ _06405_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[15]$_DFFE_PP0P_  clock_i _00638_ \atbs_core_0.spike_memory_0.n1953_o[15]\ _06404_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[16]$_DFFE_PP0P_  clock_i _00639_ \atbs_core_0.spike_memory_0.n1953_o[16]\ _06403_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[17]$_DFFE_PP0P_  clock_i _00640_ \atbs_core_0.spike_memory_0.n1953_o[17]\ _06402_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[18]$_DFFE_PP0P_  clock_i _00641_ \atbs_core_0.spike_memory_0.n1953_o[18]\ _06401_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[19]$_DFFE_PP0P_  clock_i _00642_ \atbs_core_0.spike_memory_0.n1954_o[0]\ _06400_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[1]$_DFFE_PP0P_  clock_i _00643_ \atbs_core_0.spike_memory_0.n1953_o[1]\ _06399_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[20]$_DFFE_PP0P_  clock_i _00644_ \atbs_core_0.spike_memory_0.n1954_o[1]\ _06398_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[21]$_DFFE_PP0P_  clock_i _00645_ \atbs_core_0.spike_memory_0.n1954_o[2]\ _06397_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[22]$_DFFE_PP0P_  clock_i _00646_ \atbs_core_0.spike_memory_0.n1954_o[3]\ _06396_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[23]$_DFFE_PP0P_  clock_i _00647_ \atbs_core_0.spike_memory_0.n1954_o[4]\ _06395_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[24]$_DFFE_PP0P_  clock_i _00648_ \atbs_core_0.spike_memory_0.n1954_o[5]\ _06394_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[25]$_DFFE_PP0P_  clock_i _00649_ \atbs_core_0.spike_memory_0.n1954_o[6]\ _06393_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[26]$_DFFE_PP0P_  clock_i _00650_ \atbs_core_0.spike_memory_0.n1954_o[7]\ _06392_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[27]$_DFFE_PP0P_  clock_i _00651_ \atbs_core_0.spike_memory_0.n1954_o[8]\ _06391_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[28]$_DFFE_PP0P_  clock_i _00652_ \atbs_core_0.spike_memory_0.n1954_o[9]\ _06390_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[29]$_DFFE_PP0P_  clock_i _00653_ \atbs_core_0.spike_memory_0.n1954_o[10]\ _06389_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[2]$_DFFE_PP0P_  clock_i _00654_ \atbs_core_0.spike_memory_0.n1953_o[2]\ _06388_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[30]$_DFFE_PP0P_  clock_i _00655_ \atbs_core_0.spike_memory_0.n1954_o[11]\ _06387_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[31]$_DFFE_PP0P_  clock_i _00656_ \atbs_core_0.spike_memory_0.n1954_o[12]\ _06386_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[32]$_DFFE_PP0P_  clock_i _00657_ \atbs_core_0.spike_memory_0.n1954_o[13]\ _06385_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[33]$_DFFE_PP0P_  clock_i _00658_ \atbs_core_0.spike_memory_0.n1954_o[14]\ _06384_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[34]$_DFFE_PP0P_  clock_i _00659_ \atbs_core_0.spike_memory_0.n1954_o[15]\ _06383_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[35]$_DFFE_PP0P_  clock_i _00660_ \atbs_core_0.spike_memory_0.n1954_o[16]\ _06382_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[36]$_DFFE_PP0P_  clock_i _00661_ \atbs_core_0.spike_memory_0.n1954_o[17]\ _06381_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[37]$_DFFE_PP0P_  clock_i _00662_ \atbs_core_0.spike_memory_0.n1954_o[18]\ _06380_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[38]$_DFFE_PP0P_  clock_i _00663_ \atbs_core_0.spike_memory_0.n1955_o[0]\ _06379_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[39]$_DFFE_PP0P_  clock_i _00664_ \atbs_core_0.spike_memory_0.n1955_o[1]\ _06378_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[3]$_DFFE_PP0P_  clock_i _00665_ \atbs_core_0.spike_memory_0.n1953_o[3]\ _06377_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[40]$_DFFE_PP0P_  clock_i _00666_ \atbs_core_0.spike_memory_0.n1955_o[2]\ _06376_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[41]$_DFFE_PP0P_  clock_i _00667_ \atbs_core_0.spike_memory_0.n1955_o[3]\ _06375_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[42]$_DFFE_PP0P_  clock_i _00668_ \atbs_core_0.spike_memory_0.n1955_o[4]\ _06374_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[43]$_DFFE_PP0P_  clock_i _00669_ \atbs_core_0.spike_memory_0.n1955_o[5]\ _06373_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[44]$_DFFE_PP0P_  clock_i _00670_ \atbs_core_0.spike_memory_0.n1955_o[6]\ _06372_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[45]$_DFFE_PP0P_  clock_i _00671_ \atbs_core_0.spike_memory_0.n1955_o[7]\ _06371_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[46]$_DFFE_PP0P_  clock_i _00672_ \atbs_core_0.spike_memory_0.n1955_o[8]\ _06370_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[47]$_DFFE_PP0P_  clock_i _00673_ \atbs_core_0.spike_memory_0.n1955_o[9]\ _06369_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[48]$_DFFE_PP0P_  clock_i _00674_ \atbs_core_0.spike_memory_0.n1955_o[10]\ _06368_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[49]$_DFFE_PP0P_  clock_i _00675_ \atbs_core_0.spike_memory_0.n1955_o[11]\ _06367_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[4]$_DFFE_PP0P_  clock_i _00676_ \atbs_core_0.spike_memory_0.n1953_o[4]\ _06366_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[50]$_DFFE_PP0P_  clock_i _00677_ \atbs_core_0.spike_memory_0.n1955_o[12]\ _06365_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[51]$_DFFE_PP0P_  clock_i _00678_ \atbs_core_0.spike_memory_0.n1955_o[13]\ _06364_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[52]$_DFFE_PP0P_  clock_i _00679_ \atbs_core_0.spike_memory_0.n1955_o[14]\ _06363_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[53]$_DFFE_PP0P_  clock_i _00680_ \atbs_core_0.spike_memory_0.n1955_o[15]\ _06362_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[54]$_DFFE_PP0P_  clock_i _00681_ \atbs_core_0.spike_memory_0.n1955_o[16]\ _06361_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[55]$_DFFE_PP0P_  clock_i _00682_ \atbs_core_0.spike_memory_0.n1955_o[17]\ _06360_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[56]$_DFFE_PP0P_  clock_i _00683_ \atbs_core_0.spike_memory_0.n1955_o[18]\ _06359_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[57]$_DFFE_PP0P_  clock_i _00684_ \atbs_core_0.spike_memory_0.n1971_q[57]\ _06358_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[58]$_DFFE_PP0P_  clock_i _00685_ \atbs_core_0.spike_memory_0.n1971_q[58]\ _06357_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[59]$_DFFE_PP0P_  clock_i _00686_ \atbs_core_0.spike_memory_0.n1971_q[59]\ _06356_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[5]$_DFFE_PP0P_  clock_i _00687_ \atbs_core_0.spike_memory_0.n1953_o[5]\ _06355_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[60]$_DFFE_PP0P_  clock_i _00688_ \atbs_core_0.spike_memory_0.n1971_q[60]\ _06354_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[61]$_DFFE_PP0P_  clock_i _00689_ \atbs_core_0.spike_memory_0.n1971_q[61]\ _06353_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[62]$_DFFE_PP0P_  clock_i _00690_ \atbs_core_0.spike_memory_0.n1971_q[62]\ _06352_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[63]$_DFFE_PP0P_  clock_i _00691_ \atbs_core_0.spike_memory_0.n1971_q[63]\ _06351_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[64]$_DFFE_PP0P_  clock_i _00692_ \atbs_core_0.spike_memory_0.n1971_q[64]\ _06350_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[65]$_DFFE_PP0P_  clock_i _00693_ \atbs_core_0.spike_memory_0.n1971_q[65]\ _06349_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[66]$_DFFE_PP0P_  clock_i _00694_ \atbs_core_0.spike_memory_0.n1971_q[66]\ _06348_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[67]$_DFFE_PP0P_  clock_i _00695_ \atbs_core_0.spike_memory_0.n1971_q[67]\ _06347_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[68]$_DFFE_PP0P_  clock_i _00696_ \atbs_core_0.spike_memory_0.n1971_q[68]\ _06346_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[69]$_DFFE_PP0P_  clock_i _00697_ \atbs_core_0.spike_memory_0.n1971_q[69]\ _06345_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[6]$_DFFE_PP0P_  clock_i _00698_ \atbs_core_0.spike_memory_0.n1953_o[6]\ _06344_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[70]$_DFFE_PP0P_  clock_i _00699_ \atbs_core_0.spike_memory_0.n1971_q[70]\ _06343_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[71]$_DFFE_PP0P_  clock_i _00700_ \atbs_core_0.spike_memory_0.n1971_q[71]\ _06342_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[72]$_DFFE_PP0P_  clock_i _00701_ \atbs_core_0.spike_memory_0.n1971_q[72]\ _06341_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[73]$_DFFE_PP0P_  clock_i _00702_ \atbs_core_0.spike_memory_0.n1971_q[73]\ _06340_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[74]$_DFFE_PP0P_  clock_i _00703_ \atbs_core_0.spike_memory_0.n1971_q[74]\ _06339_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[75]$_DFFE_PP0P_  clock_i _00704_ \atbs_core_0.spike_memory_0.n1971_q[75]\ _06338_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[7]$_DFFE_PP0P_  clock_i _00705_ \atbs_core_0.spike_memory_0.n1953_o[7]\ _06337_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[8]$_DFFE_PP0P_  clock_i _00706_ \atbs_core_0.spike_memory_0.n1953_o[8]\ _06336_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1971_q[9]$_DFFE_PP0P_  clock_i _00707_ \atbs_core_0.spike_memory_0.n1953_o[9]\ _06335_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1972_q[0]$_DFFE_PP0P_  clock_i _00708_ \atbs_core_0.spike_memory_0.head[0]\ \atbs_core_0.spike_memory_0.n1901_o[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1972_q[1]$_DFFE_PP0P_  clock_i _00709_ \atbs_core_0.spike_memory_0.head[1]\ _06334_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1973_q[0]$_DFFE_PP0P_  clock_i _00710_ \atbs_core_0.spike_memory_0.n1973_q[0]\ \atbs_core_0.spike_memory_0.n1916_o[0]\ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1973_q[1]$_DFFE_PP0P_  clock_i _00711_ \atbs_core_0.spike_memory_0.n1973_q[1]\ _06333_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1974_q$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1899_o\ \atbs_core_0.spike_memory_0.n1974_q\ _06332_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[0]$_DFFE_PP0P_  clock_i _00712_ \atbs_core_0.spike_memory_0.a_data[0]\ _06331_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[10]$_DFFE_PP0P_  clock_i _00713_ \atbs_core_0.spike_memory_0.a_data[10]\ _06330_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[11]$_DFFE_PP0P_  clock_i _00714_ \atbs_core_0.spike_memory_0.a_data[11]\ _06329_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[12]$_DFFE_PP0P_  clock_i _00715_ \atbs_core_0.spike_memory_0.a_data[12]\ _06328_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[13]$_DFFE_PP0P_  clock_i _00716_ \atbs_core_0.spike_memory_0.a_data[13]\ _06327_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[14]$_DFFE_PP0P_  clock_i _00717_ \atbs_core_0.spike_memory_0.a_data[14]\ _06326_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[15]$_DFFE_PP0P_  clock_i _00718_ \atbs_core_0.spike_memory_0.a_data[15]\ _06325_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[16]$_DFFE_PP0P_  clock_i _00719_ \atbs_core_0.spike_memory_0.a_data[16]\ _06324_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[17]$_DFFE_PP0P_  clock_i _00720_ \atbs_core_0.spike_memory_0.a_data[17]\ _06323_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[18]$_DFFE_PP0P_  clock_i _00721_ \atbs_core_0.spike_memory_0.a_data[18]\ _06322_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[1]$_DFFE_PP0P_  clock_i _00722_ \atbs_core_0.spike_memory_0.a_data[1]\ _06321_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[2]$_DFFE_PP0P_  clock_i _00723_ \atbs_core_0.spike_memory_0.a_data[2]\ _06320_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[3]$_DFFE_PP0P_  clock_i _00724_ \atbs_core_0.spike_memory_0.a_data[3]\ _06319_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[4]$_DFFE_PP0P_  clock_i _00725_ \atbs_core_0.spike_memory_0.a_data[4]\ _06318_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[5]$_DFFE_PP0P_  clock_i _00726_ \atbs_core_0.spike_memory_0.a_data[5]\ _06317_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[6]$_DFFE_PP0P_  clock_i _00727_ \atbs_core_0.spike_memory_0.a_data[6]\ _06316_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[7]$_DFFE_PP0P_  clock_i _00728_ \atbs_core_0.spike_memory_0.a_data[7]\ _06315_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[8]$_DFFE_PP0P_  clock_i _00729_ \atbs_core_0.spike_memory_0.a_data[8]\ _06314_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1975_q[9]$_DFFE_PP0P_  clock_i _00730_ \atbs_core_0.spike_memory_0.a_data[9]\ _06313_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[0]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[0]\ \atbs_core_0.b_data[0]\ _06312_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[10]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[10]\ \atbs_core_0.b_data[10]\ _06311_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[11]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[11]\ \atbs_core_0.b_data[11]\ _06310_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[12]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[12]\ \atbs_core_0.b_data[12]\ _06309_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[13]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[13]\ \atbs_core_0.b_data[13]\ _06308_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[14]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[14]\ \atbs_core_0.b_data[14]\ _06307_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[15]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[15]\ \atbs_core_0.b_data[15]\ _06306_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[16]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[16]\ \atbs_core_0.b_data[16]\ _06305_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[17]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[17]\ \atbs_core_0.b_data[17]\ _06304_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[18]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[18]\ \atbs_core_0.b_data[18]\ _06303_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[1]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[1]\ \atbs_core_0.b_data[1]\ _06302_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[2]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[2]\ \atbs_core_0.b_data[2]\ _06301_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[3]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[3]\ \atbs_core_0.b_data[3]\ _06300_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[4]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[4]\ \atbs_core_0.b_data[4]\ _06299_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[5]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[5]\ \atbs_core_0.b_data[5]\ _06298_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[6]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[6]\ \atbs_core_0.b_data[6]\ _06297_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[7]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[7]\ \atbs_core_0.b_data[7]\ _06296_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[8]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[8]\ \atbs_core_0.b_data[8]\ _06295_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1976_q[9]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1985_o[9]\ \atbs_core_0.b_data[9]\ _06294_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1977_q[0]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1914_o\ \atbs_core_0.spike_memory_0.n1968_o\ _06293_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1977_q[1]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1968_o\ \atbs_core_0.spike_memory_0.n1966_o\ _06292_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1977_q[2]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1966_o\ \atbs_core_0.spike_memory_0.n1964_o\ _06291_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1977_q[3]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n1964_o\ \atbs_core_0.memory2uart_0.read_strb_i\ _06290_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1979_q[0]$_DFFE_PP0P_  clock_i _00731_ \atbs_core_0.spike_memory_0.n1926_o\ _06289_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1979_q[1]$_DFFE_PP0P_  clock_i _00732_ \atbs_core_0.spike_memory_0.n1925_o\ _06288_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n1979_q[2]$_DFFE_PP0P_  clock_i _00733_ \atbs_core_0.spike_memory_0.n1912_o\ _06935_ _00119_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_0.n1095_q[0]$_DFF_PN0_  clock_i _06940_ \atbs_core_0.sync_chain_0.n1088_o\ _06936_ reset_n_i VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_0.n1095_q[1]$_DFF_PN0_  clock_i \atbs_core_0.sync_chain_0.n1088_o\ \atbs_core_0.n31_o\ _06287_ reset_n_i VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1187_q[0]$_DFF_PP0_  clock_i comp_upper_i \atbs_core_0.sync_chain_1.buf[0]\ _06286_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1187_q[1]$_DFF_PP0_  clock_i comp_lower_i \atbs_core_0.sync_chain_1.buf[1]\ _06285_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1187_q[2]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_1.buf[0]\ \atbs_core_0.comp_upper_sync\ _06284_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1187_q[3]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_1.buf[1]\ \atbs_core_0.comp_lower_sync\ _06283_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_2.n1095_q[0]$_DFF_PP0_  clock_i trigger_start_sampling_i \atbs_core_0.sync_chain_2.n1088_o\ _06282_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_2.n1095_q[1]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_2.n1088_o\ \atbs_core_0.n37_o\ _06281_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[0]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[0]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[0]\ _00061_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[10]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[10]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[10]\ _00017_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[11]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[11]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[11]\ _00016_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[12]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[12]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[12]\ _00015_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[13]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[13]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[13]\ _00014_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[14]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[14]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[14]\ _00013_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[15]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[15]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[15]\ _00012_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[16]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[16]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[16]\ _00021_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[17]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[17]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[17]\ _00020_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[1]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[1]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[1]\ _00062_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[2]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[2]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[2]\ _00063_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[3]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[3]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[3]\ _00064_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[4]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[4]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[4]\ _00065_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[5]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[5]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[5]\ _00066_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[6]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[6]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[6]\ _00011_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[7]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[7]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[7]\ _00010_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[8]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[8]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[8]\ _00019_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1818_q[9]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1813_o[9]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[9]\ _00018_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n1819_q$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n1809_o\ \atbs_core_0.adaptive_ctrl_0.n1308_o\ _00052_ _00122_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2883_q[0]$_DFFE_PP0P_  clock_i _00734_ \atbs_core_0.uart_0.uart_rx_0.n2897_o\ _00007_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2883_q[1]$_DFFE_PP0P_  clock_i _00735_ \atbs_core_0.uart_0.uart_rx_0.n2891_o\ _06280_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2883_q[2]$_DFFE_PP0P_  clock_i _00736_ \atbs_core_0.uart_0.uart_rx_0.n2889_o\ _06279_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[0]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[0]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[0]\ _06278_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[1]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[1]\ _06277_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[2]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[2]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[2]\ _06276_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[3]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[3]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ _06275_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[4]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[4]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[4]\ _06274_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[5]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[5]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[5]\ _06273_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[6]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[6]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[6]\ _06272_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[7]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[7]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ _06271_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2884_q[8]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2836_o[8]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ _00006_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[0]$_DFFE_PP0P_  clock_i _00737_ \atbs_core_0.uart_0.uart_rx_0.n2907_o\ _06270_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[1]$_DFFE_PP0P_  clock_i _00738_ \atbs_core_0.uart_0.uart_rx_0.n2909_o\ _06269_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[2]$_DFFE_PP0P_  clock_i _00739_ \atbs_core_0.uart_0.uart_rx_0.n2911_o\ _06268_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[3]$_DFFE_PP0P_  clock_i _00740_ \atbs_core_0.uart_0.uart_rx_0.n2913_o\ _06267_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[4]$_DFFE_PP0P_  clock_i _00741_ \atbs_core_0.uart_0.uart_rx_0.n2915_o\ _06266_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[5]$_DFFE_PP0P_  clock_i _00742_ \atbs_core_0.uart_0.uart_rx_0.n2917_o\ _06265_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[6]$_DFFE_PP0P_  clock_i _00743_ \atbs_core_0.uart_0.uart_rx_0.n2919_o\ _06264_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2885_q[7]$_DFFE_PP0P_  clock_i _00744_ \atbs_core_0.uart_0.uart_rx_0.n2921_o\ _06263_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2886_q$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n2880_o\ \atbs_core_0.uart_0.rx_data_strb_o\ _06262_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2887_q[0]$_DFF_PP1_  clock_i _00123_ _06938_ \atbs_core_0.uart_0.uart_rx_0.n2834_o\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2887_q[1]$_DFF_PP0_  clock_i _00000_ \atbs_core_0.uart_0.uart_rx_0.n2819_o\ _06261_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2887_q[2]$_DFF_PP0_  clock_i _00001_ \atbs_core_0.uart_0.uart_rx_0.n2848_o\ _06260_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n2887_q[3]$_DFF_PP0_  clock_i _00002_ \atbs_core_0.uart_0.uart_rx_0.n2873_o\ _06259_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2779_q$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2776_o\ \atbs_core_0.memory2uart_0.tx_strb_i\ \atbs_core_0.spike_memory_0.n1928_o[0]\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2780_q[0]$_DFFE_PP0P_  clock_i _00745_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[0]\ _06258_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2780_q[1]$_DFFE_PP0P_  clock_i _00746_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[1]\ _06257_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2780_q[2]$_DFFE_PP0P_  clock_i _00747_ \atbs_core_0.uart_0.uart_tx_0.n2780_q[2]\ _00060_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[0]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[0]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[0]\ _06256_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[1]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[1]\ _06255_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[2]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[2]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[2]\ _06254_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[3]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[3]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[3]\ _06253_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[4]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[4]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[4]\ _06252_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[5]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[5]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[5]\ _06251_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[6]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[6]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ _06250_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[7]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[7]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[7]\ _06249_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2781_q[8]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2712_o[8]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[8]\ _06248_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2782_q[0]$_DFF_PP1_  clock_i _00124_ _06939_ \atbs_core_0.uart_0.uart_tx_0.n2721_o\ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2782_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n2766_o[2]\ \atbs_core_0.uart_0.uart_tx_0.n2758_o\ _00022_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2782_q[2]$_DFF_PP0_  clock_i _00003_ \atbs_core_0.uart_0.uart_tx_0.n2735_o\ _06247_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2782_q[3]$_DFF_PP0_  clock_i _00004_ \atbs_core_0.uart_0.uart_tx_0.n2730_o\ _06246_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n2782_q[4]$_DFF_PP0_  clock_i _00005_ \atbs_core_0.uart_0.uart_tx_0.n2699_o\ _06245_ _00120_ VPWR 
+ VGND
+ sg13g2_dfrbp_1

.ends
.end
