*SPICE netlist created from verilog structural netlist module atbs_core_fixed_window_board by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

.subckt atbs_core_fixed_window_board VPWR VGND adaptive_mode_i bio_amp_en_o clock_i comp_lower_i comp_upper_i
+ control_mode_i dac_lower_o[0] dac_lower_o[1] dac_lower_o[2] dac_lower_o[3] dac_upper_o[0] dac_upper_o[1] dac_upper_o[2]
+ dac_upper_o[3] enable_i idle_led_o overflow_led_o phi_bias_1_o phi_bias_2_o phi_cmfb_1_o phi_cmfb_2_o
+ phi_comp_o phi_dac_lower_o phi_dac_upper_o phi_res_1_o phi_res_2_o phi_vcm_generator_1_o phi_vcm_generator_2_o reset_n_i
+ select_cap_o[0] select_cap_o[1] select_cap_o[2] select_spdt_o select_tbs_delta_steps_i signal_select_in_i spike_o trigger_start_mode_i
+ trigger_start_sampling_i uart_rx_i uart_tx_o underflow_led_o 

X_14578_ \atbs_core_0.enable_read\ VPWR VGND _07516_ sg13g2_inv_1
X_14579_ \atbs_core_0.spike_memory_0.head[3]\ VPWR VGND _07517_ sg13g2_buf_1
X_14580_ \atbs_core_0.spike_memory_0.n2438_q[3]\ VPWR VGND _07518_ sg13g2_buf_1
X_14581_ \atbs_core_0.spike_memory_0.n2438_q[2]\ VPWR VGND _07519_ sg13g2_buf_1
X_14582_ \atbs_core_0.spike_memory_0.head[2]\ VPWR VGND _07520_ sg13g2_buf_1
X_14583_ _07519_ _07520_ VPWR VGND _07521_ sg13g2_nor2b_1
X_14584_ \atbs_core_0.spike_memory_0.n2438_q[1]\ VPWR VGND _07522_ sg13g2_buf_1
X_14585_ \atbs_core_0.spike_memory_0.head[1]\ VPWR VGND _07523_ sg13g2_buf_1
X_14586_ _07522_ _07523_ VPWR VGND _07524_ sg13g2_nand2b_1
X_14587_ \atbs_core_0.spike_memory_0.head[0]\ VPWR VGND _07525_ sg13g2_buf_1
X_14588_ \atbs_core_0.spike_memory_0.n2438_q[0]\ VPWR VGND _07526_ sg13g2_buf_2
X_14589_ _07525_ _07526_ VPWR VGND _07527_ sg13g2_nor2b_1
X_14590_ _07527_ VPWR VGND _07528_ sg13g2_buf_1
X_14591_ _07523_ _07522_ VPWR VGND _07529_ sg13g2_nor2b_1
X_14592_ _07524_ _07528_ _07529_ VPWR VGND _07530_ sg13g2_a21oi_1
X_14593_ _07520_ _07519_ VPWR VGND _07531_ sg13g2_nand2b_1
X_14594_ _07521_ _07530_ _07531_ VPWR VGND _07532_ sg13g2_o21ai_1
X_14595_ _07532_ VPWR VGND _07533_ sg13g2_buf_1
X_14596_ _07518_ _07533_ VPWR VGND _07534_ sg13g2_nand2_1
X_14597_ _07518_ _07533_ VPWR VGND _07535_ sg13g2_nor2_1
X_14598_ _07517_ _07534_ _07535_ VPWR VGND _07536_ sg13g2_a21oi_1
X_14599_ \atbs_core_0.spike_memory_0.head[4]\ VPWR VGND _07537_ sg13g2_buf_1
X_14600_ \atbs_core_0.spike_memory_0.n2438_q[4]\ VPWR VGND _07538_ sg13g2_buf_1
X_14601_ _07537_ _07538_ VPWR VGND _07539_ sg13g2_xor2_1
X_14602_ _07536_ _07539_ VPWR VGND _07540_ sg13g2_xnor2_1
X_14603_ _07540_ VPWR VGND _07541_ sg13g2_buf_1
X_14604_ \atbs_core_0.spike_memory_0.head[5]\ \atbs_core_0.spike_memory_0.n2438_q[5]\ VPWR VGND _07542_ sg13g2_xor2_1
X_14605_ _07538_ _07536_ VPWR VGND _07543_ sg13g2_nand2_1
X_14606_ _07538_ _07536_ VPWR VGND _07544_ sg13g2_nor2_1
X_14607_ _07537_ _07543_ _07544_ VPWR VGND _07545_ sg13g2_a21oi_1
X_14608_ _07542_ _07545_ VPWR VGND _07546_ sg13g2_xnor2_1
X_14609_ _07546_ VPWR VGND _07547_ sg13g2_buf_1
X_14610_ _07541_ _07547_ VPWR VGND _07548_ sg13g2_nand2_1
X_14611_ _07548_ VPWR VGND _07549_ sg13g2_buf_2
X_14612_ _07521_ _07531_ VPWR VGND _07550_ sg13g2_nor2b_1
X_14613_ _07530_ _07550_ VPWR VGND _07551_ sg13g2_xnor2_1
X_14614_ _07551_ VPWR VGND _07552_ sg13g2_buf_1
X_14615_ _07517_ _07518_ VPWR VGND _07553_ sg13g2_xnor2_1
X_14616_ _07533_ _07553_ VPWR VGND _07554_ sg13g2_xor2_1
X_14617_ _07554_ VPWR VGND _07555_ sg13g2_buf_1
X_14618_ _07552_ _07555_ VPWR VGND _07556_ sg13g2_nand2_1
X_14619_ _07523_ _07522_ VPWR VGND _07557_ sg13g2_xnor2_1
X_14620_ _07557_ VPWR VGND _07558_ sg13g2_buf_1
X_14621_ _07526_ _07525_ VPWR VGND _07559_ sg13g2_nor2b_1
X_14622_ _07559_ VPWR VGND _07560_ sg13g2_buf_1
X_14623_ _07528_ _07560_ VPWR VGND _07561_ sg13g2_nor2_1
X_14624_ _07558_ _07561_ VPWR VGND _07562_ sg13g2_nand2_1
X_14625_ _07562_ VPWR VGND _07563_ sg13g2_buf_1
X_14626_ _07549_ _07556_ _07563_ VPWR VGND _07564_ sg13g2_nor3_1
X_14627_ _07516_ \atbs_core_0.spike_memory_0.n2317_o\ _07564_ VPWR VGND _07565_ sg13g2_nor3_1
X_14628_ _07565_ VPWR VGND \atbs_core_0.spike_memory_0.n2319_o\ sg13g2_buf_2
X_14629_ \atbs_core_0.spike_detector_0.n1595_q\ \atbs_core_0.spike_detector_0.lower_is_changing\ VPWR VGND _07566_ sg13g2_nor2_1
X_14630_ _07566_ VPWR VGND \atbs_core_0.spike_detector_0.n1583_o\ sg13g2_inv_1
X_14631_ \atbs_core_0.uart_0.uart_rx_0.n3413_o\ VPWR VGND _07567_ sg13g2_buf_1
X_14632_ _07567_ VPWR VGND _07568_ sg13g2_inv_1
X_14633_ \atbs_core_0.baudrate_adj_uart[7]\ VPWR VGND _07569_ sg13g2_buf_1
X_14634_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ VPWR VGND _07570_ sg13g2_inv_1
X_14635_ _07569_ _07570_ VPWR VGND _07571_ sg13g2_nor2_1
X_14636_ _07569_ _07570_ VPWR VGND _07572_ sg13g2_nand2_1
X_14637_ _07571_ _07572_ VPWR VGND _07573_ sg13g2_nor2b_1
X_14638_ \atbs_core_0.baudrate_adj_uart[6]\ VPWR VGND _07574_ sg13g2_buf_1
X_14639_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[6]\ VPWR VGND _07575_ sg13g2_buf_1
X_14640_ _07574_ _07575_ VPWR VGND _07576_ sg13g2_xnor2_1
X_14641_ \atbs_core_0.baudrate_adj_uart[2]\ VPWR VGND _07577_ sg13g2_buf_1
X_14642_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[2]\ VPWR VGND _07578_ sg13g2_buf_1
X_14643_ _07577_ _07578_ VPWR VGND _07579_ sg13g2_xnor2_1
X_14644_ \atbs_core_0.baudrate_adj_uart[5]\ VPWR VGND _07580_ sg13g2_buf_1
X_14645_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[5]\ VPWR VGND _07581_ sg13g2_buf_1
X_14646_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ VPWR VGND _07582_ sg13g2_buf_1
X_14647_ _07580_ _07581_ _07582_ VPWR VGND _07583_ sg13g2_nand3_1
X_14648_ _07580_ _07581_ _07582_ VPWR VGND _07584_ sg13g2_or3_1
X_14649_ \atbs_core_0.baudrate_adj_uart[1]\ VPWR VGND _07585_ sg13g2_buf_1
X_14650_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[1]\ VPWR VGND _07586_ sg13g2_buf_1
X_14651_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ VPWR VGND _07587_ sg13g2_buf_1
X_14652_ _07585_ _07586_ _07587_ VPWR VGND _07588_ sg13g2_nand3_1
X_14653_ _07585_ _07586_ _07587_ VPWR VGND _07589_ sg13g2_or3_1
X_14654_ \atbs_core_0.baudrate_adj_uart[4]\ VPWR VGND _07590_ sg13g2_buf_1
X_14655_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[4]\ VPWR VGND _07591_ sg13g2_buf_1
X_14656_ _07590_ _07591_ VPWR VGND _07592_ sg13g2_nand2b_1
X_14657_ _07591_ _07590_ VPWR VGND _07593_ sg13g2_nand2b_1
X_14658_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[0]\ VPWR VGND _07594_ sg13g2_buf_1
X_14659_ \atbs_core_0.baudrate_adj_uart[0]\ VPWR VGND _07595_ sg13g2_buf_1
X_14660_ _07594_ _07595_ VPWR VGND _07596_ sg13g2_nand2b_1
X_14661_ _07595_ _07594_ VPWR VGND _07597_ sg13g2_nand2b_1
X_14662_ _07592_ _07593_ _07596_ _07597_ VPWR VGND 
+ _07598_
+ sg13g2_nand4_1
X_14663_ _07583_ _07584_ _07588_ _07589_ _07598_ VPWR 
+ VGND
+ _07599_ sg13g2_a221oi_1
X_14664_ _07573_ _07576_ _07579_ _07599_ VPWR VGND 
+ _07600_
+ sg13g2_nand4_1
X_14665_ _07600_ VPWR VGND _07601_ sg13g2_buf_1
X_14666_ \atbs_core_0.uart_0.uart_rx_0.n3456_o\ VPWR VGND _07602_ sg13g2_buf_1
X_14667_ \atbs_core_0.uart_0.uart_rx_0.n3454_o\ VPWR VGND _07603_ sg13g2_buf_1
X_14668_ _07602_ _07603_ VPWR VGND _07604_ sg13g2_nand2_1
X_14669_ \atbs_core_0.uart_0.uart_rx_0.n3462_o\ VPWR VGND _07605_ sg13g2_buf_1
X_14670_ _07601_ VPWR VGND _07606_ sg13g2_inv_1
X_14671_ _07605_ _07606_ VPWR VGND _07607_ sg13g2_nand2_1
X_14672_ \atbs_core_0.uart_0.uart_rx_0.n3384_o\ VPWR VGND _07608_ sg13g2_buf_1
X_14673_ _07604_ _07607_ _07608_ VPWR VGND _07609_ sg13g2_o21ai_1
X_14674_ _07568_ _07601_ _07609_ VPWR VGND _00000_ sg13g2_o21ai_1
X_14675_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[5]\ VPWR VGND _07610_ sg13g2_buf_1
X_14676_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[8]\ VPWR VGND _07611_ sg13g2_buf_1
X_14677_ _07610_ _07611_ VPWR VGND _07612_ sg13g2_or2_1
X_14678_ _07580_ _07610_ _07611_ VPWR VGND _07613_ sg13g2_nand3_1
X_14679_ _07580_ _07612_ _07613_ VPWR VGND _07614_ sg13g2_o21ai_1
X_14680_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[0]\ VPWR VGND _07615_ sg13g2_buf_1
X_14681_ _07595_ _07615_ VPWR VGND _07616_ sg13g2_nand2b_1
X_14682_ _07574_ VPWR VGND _07617_ sg13g2_inv_1
X_14683_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ VPWR VGND _07618_ sg13g2_buf_1
X_14684_ _07617_ _07618_ VPWR VGND _07619_ sg13g2_nand2_1
X_14685_ _07618_ _07574_ VPWR VGND _07620_ sg13g2_nand2b_1
X_14686_ _07614_ _07616_ _07619_ _07620_ VPWR VGND 
+ _07621_
+ sg13g2_nand4_1
X_14687_ _07585_ VPWR VGND _07622_ sg13g2_inv_1
X_14688_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[1]\ VPWR VGND _07623_ sg13g2_buf_1
X_14689_ _07615_ VPWR VGND _07624_ sg13g2_inv_1
X_14690_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[2]\ VPWR VGND _07625_ sg13g2_buf_1
X_14691_ _07577_ _07625_ VPWR VGND _07626_ sg13g2_xor2_1
X_14692_ _07595_ _07624_ _07623_ _07622_ _07626_ VPWR 
+ VGND
+ _07627_ sg13g2_a221oi_1
X_14693_ _07622_ _07623_ _07627_ VPWR VGND _07628_ sg13g2_o21ai_1
X_14694_ _07569_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[7]\ VPWR VGND _07629_ sg13g2_xnor2_1
X_14695_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[3]\ VPWR VGND _07630_ sg13g2_buf_1
X_14696_ _07585_ _07630_ VPWR VGND _07631_ sg13g2_xnor2_1
X_14697_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[4]\ VPWR VGND _07632_ sg13g2_buf_1
X_14698_ _07590_ _07632_ VPWR VGND _07633_ sg13g2_nand2b_1
X_14699_ _07632_ _07590_ VPWR VGND _07634_ sg13g2_nand2b_1
X_14700_ _07629_ _07631_ _07633_ _07634_ VPWR VGND 
+ _07635_
+ sg13g2_nand4_1
X_14701_ _07621_ _07628_ _07635_ VPWR VGND _07636_ sg13g2_nor3_1
X_14702_ _07636_ VPWR VGND _07637_ sg13g2_buf_1
X_14703_ \atbs_core_0.uart_0.uart_tx_0.n3286_o\ VPWR VGND _07638_ sg13g2_buf_1
X_14704_ _00062_ VPWR VGND _07639_ sg13g2_inv_1
X_14705_ \atbs_core_0.uart_0.uart_tx_0.n3295_o\ VPWR VGND _07640_ sg13g2_buf_1
X_14706_ _07638_ _07639_ _07640_ VPWR VGND _07641_ sg13g2_a21oi_1
X_14707_ _07637_ _07641_ VPWR VGND _00004_ sg13g2_nor2_1
X_14708_ \atbs_core_0.uart_0.uart_tx_0.n3300_o\ VPWR VGND _07642_ sg13g2_buf_1
X_14709_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[1]\ VPWR VGND _07643_ sg13g2_buf_1
X_14710_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[0]\ VPWR VGND _07644_ sg13g2_buf_1
X_14711_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[2]\ VPWR VGND _07645_ sg13g2_buf_1
X_14712_ _07643_ _07644_ _07645_ _07637_ VPWR VGND 
+ _07646_
+ sg13g2_nand4_1
X_14713_ \atbs_core_0.uart_0.uart_tx_0.n3264_o\ VPWR VGND _07647_ sg13g2_buf_1
X_14714_ _07642_ _07637_ _07646_ _07647_ VPWR VGND 
+ _07648_
+ sg13g2_a22oi_1
X_14715_ _07648_ VPWR VGND _00005_ sg13g2_inv_1
X_14716_ \atbs_core_0.uart_0.uart_tx_0.n3323_o\ VPWR VGND _07649_ sg13g2_buf_1
X_14717_ _07638_ _07649_ \atbs_core_0.memory2uart_0.n2605_q\ VPWR VGND _07650_ sg13g2_o21ai_1
X_14718_ _07640_ _07650_ VPWR VGND _07651_ sg13g2_nor2b_1
X_14719_ _07642_ _07637_ VPWR VGND _07652_ sg13g2_nor2_1
X_14720_ _07637_ _07651_ _07652_ VPWR VGND _00003_ sg13g2_a21oi_1
X_14721_ \atbs_core_0.control_mode_debounced\ VPWR VGND _07653_ sg13g2_buf_16
X_14722_ _07653_ \atbs_core_0.debouncer_4.debounced\ VPWR VGND _07654_ sg13g2_nor2b_1
X_14723_ _07653_ \atbs_core_0.enable_analog_uart\ _07654_ VPWR VGND _07655_ sg13g2_a21oi_1
X_14724_ _07655_ VPWR VGND _07656_ sg13g2_inv_1
X_14725_ _07656_ VPWR VGND _07657_ sg13g2_buf_1
X_14726_ _07657_ VPWR VGND _07658_ sg13g2_buf_1
X_14727_ _07658_ VPWR VGND bio_amp_en_o sg13g2_buf_1
X_14728_ _07608_ _07602_ _07603_ VPWR VGND _07659_ sg13g2_nand3_1
X_14729_ \atbs_core_0.uart_0.uart_rx_0.n3438_o\ VPWR VGND _07660_ sg13g2_buf_1
X_14730_ _07594_ _07578_ VPWR VGND _07661_ sg13g2_or2_1
X_14731_ _07585_ _07594_ _07578_ VPWR VGND _07662_ sg13g2_nand3_1
X_14732_ _07585_ _07661_ _07662_ VPWR VGND _07663_ sg13g2_o21ai_1
X_14733_ _07575_ _07569_ VPWR VGND _07664_ sg13g2_xnor2_1
X_14734_ _00057_ _07663_ _07664_ VPWR VGND _07665_ sg13g2_nand3_1
X_14735_ _07591_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ VPWR VGND _07666_ sg13g2_or2_1
X_14736_ _07591_ _07580_ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ VPWR VGND _07667_ sg13g2_nand3_1
X_14737_ _07580_ _07666_ _07667_ VPWR VGND _07668_ sg13g2_o21ai_1
X_14738_ _07586_ _07577_ VPWR VGND _07669_ sg13g2_xor2_1
X_14739_ _07587_ _07590_ VPWR VGND _07670_ sg13g2_xor2_1
X_14740_ _07581_ _07574_ VPWR VGND _07671_ sg13g2_xor2_1
X_14741_ _07669_ _07670_ _07671_ VPWR VGND _07672_ sg13g2_nor3_1
X_14742_ _07665_ _07668_ _07672_ VPWR VGND _07673_ sg13g2_nand3b_1
X_14743_ _07660_ _07673_ VPWR VGND _07674_ sg13g2_nand2_1
X_14744_ _07607_ _07659_ _07674_ VPWR VGND _00002_ sg13g2_o21ai_1
X_14745_ \atbs_core_0.uart_0.uart_rx_0.n3399_o\ VPWR VGND _07675_ sg13g2_buf_1
X_14746_ uart_rx_i VPWR VGND _07676_ sg13g2_inv_1
X_14747_ _07675_ _07676_ _07601_ _07567_ VPWR VGND 
+ _07677_
+ sg13g2_a22oi_1
X_14748_ _07677_ VPWR VGND _00001_ sg13g2_inv_1
X_14749_ \atbs_core_0.dac_control_0.n1833_o\ VPWR VGND _07678_ sg13g2_buf_1
X_14750_ _07678_ VPWR VGND _07679_ sg13g2_buf_1
X_14751_ _07655_ VPWR VGND _07680_ sg13g2_buf_1
X_14752_ \atbs_core_0.n1412_q[2]\ VPWR VGND _07681_ sg13g2_buf_1
X_14753_ _07681_ VPWR VGND _07682_ sg13g2_inv_1
X_14754_ _07682_ _00056_ VPWR VGND _07683_ sg13g2_nand2_1
X_14755_ _07683_ VPWR VGND _07684_ sg13g2_buf_1
X_14756_ \atbs_core_0.n1412_q[1]\ VPWR VGND _07685_ sg13g2_buf_1
X_14757_ \atbs_core_0.n1412_q[0]\ _07685_ VPWR VGND _07686_ sg13g2_nand2b_1
X_14758_ \atbs_core_0.main_counter_value[8]\ VPWR VGND _07687_ sg13g2_buf_1
X_14759_ \atbs_core_0.main_counter_value[11]\ VPWR VGND _07688_ sg13g2_buf_1
X_14760_ \atbs_core_0.main_counter_value[15]\ VPWR VGND _07689_ sg13g2_buf_1
X_14761_ _07687_ _07688_ _07689_ \atbs_core_0.main_counter_value[14]\ VPWR VGND 
+ _07690_
+ sg13g2_nor4_1
X_14762_ \atbs_core_0.main_counter_value[9]\ _07690_ VPWR VGND _07691_ sg13g2_nor2b_1
X_14763_ \atbs_core_0.main_counter_value[12]\ VPWR VGND _07692_ sg13g2_buf_1
X_14764_ \atbs_core_0.main_counter_value[10]\ \atbs_core_0.main_counter_value[13]\ _07692_ VPWR VGND _07693_ sg13g2_nor3_1
X_14765_ \atbs_core_0.main_counter_value[3]\ _07691_ _07693_ VPWR VGND _07694_ sg13g2_nand3_1
X_14766_ \atbs_core_0.main_counter_value[18]\ VPWR VGND _07695_ sg13g2_buf_1
X_14767_ _07695_ \atbs_core_0.main_counter_value[19]\ VPWR VGND _07696_ sg13g2_nor2_1
X_14768_ \atbs_core_0.main_counter_value[5]\ VPWR VGND _07697_ sg13g2_buf_1
X_14769_ \atbs_core_0.main_counter_value[4]\ VPWR VGND _07698_ sg13g2_buf_1
X_14770_ _07697_ _07698_ \atbs_core_0.main_counter_value[6]\ \atbs_core_0.main_counter_value[7]\ VPWR VGND 
+ _07699_
+ sg13g2_nor4_1
X_14771_ \atbs_core_0.main_counter_value[0]\ VPWR VGND _07700_ sg13g2_buf_1
X_14772_ \atbs_core_0.main_counter_value[1]\ VPWR VGND _07701_ sg13g2_buf_1
X_14773_ _07700_ _07701_ \atbs_core_0.main_counter_value[2]\ VPWR VGND _07702_ sg13g2_nor3_1
X_14774_ _07696_ _07699_ _07702_ VPWR VGND _07703_ sg13g2_nand3_1
X_14775_ \atbs_core_0.main_counter_value[17]\ VPWR VGND _07704_ sg13g2_buf_1
X_14776_ \atbs_core_0.main_counter_value[16]\ VPWR VGND _07705_ sg13g2_buf_1
X_14777_ _07704_ _07705_ VPWR VGND _07706_ sg13g2_nor2b_1
X_14778_ _07703_ _07706_ VPWR VGND _07707_ sg13g2_nand2b_1
X_14779_ _07684_ _07686_ _07694_ _07707_ VPWR VGND 
+ _07708_
+ sg13g2_nor4_1
X_14780_ _07708_ VPWR VGND _07709_ sg13g2_buf_1
X_14781_ \atbs_core_0.adaptive_mode_debounced\ VPWR VGND _07710_ sg13g2_buf_4
X_14782_ _07710_ \atbs_core_0.adaptive_mode_uart\ _07653_ VPWR VGND _07711_ sg13g2_mux2_2
X_14783_ _07711_ VPWR VGND _07712_ sg13g2_buf_8
X_14784_ _07712_ VPWR VGND _07713_ sg13g2_buf_2
X_14785_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ VPWR VGND _07714_ sg13g2_inv_1
X_14786_ \atbs_core_0.adaptive_ctrl_0.adapt_on_overflow\ VPWR VGND _07715_ sg13g2_buf_2
X_14787_ \atbs_core_0.spike_detector_0.lock_detection\ VPWR VGND _07716_ sg13g2_buf_1
X_14788_ \atbs_core_0.detection_en\ VPWR VGND _07717_ sg13g2_inv_1
X_14789_ _07716_ _07717_ VPWR VGND _07718_ sg13g2_nor2_1
X_14790_ \atbs_core_0.adaptive_ctrl_0.n1705_o[5]\ VPWR VGND _07719_ sg13g2_buf_2
X_14791_ \atbs_core_0.adaptive_ctrl_0.n1705_o[4]\ VPWR VGND _07720_ sg13g2_buf_2
X_14792_ \atbs_core_0.adaptive_ctrl_0.n1705_o[6]\ VPWR VGND _07721_ sg13g2_buf_2
X_14793_ \atbs_core_0.adaptive_ctrl_0.n1785_q[7]\ VPWR VGND _07722_ sg13g2_buf_2
X_14794_ _07719_ _07720_ _07721_ _07722_ VPWR VGND 
+ _07723_
+ sg13g2_nor4_2
X_14795_ \atbs_core_0.adaptive_ctrl_0.n1705_o[1]\ VPWR VGND _07724_ sg13g2_buf_2
X_14796_ \atbs_core_0.adaptive_ctrl_0.n1705_o[0]\ VPWR VGND _07725_ sg13g2_buf_2
X_14797_ _07724_ _07725_ VPWR VGND _07726_ sg13g2_nor2_2
X_14798_ \atbs_core_0.adaptive_ctrl_0.n1705_o[3]\ VPWR VGND _07727_ sg13g2_buf_1
X_14799_ \atbs_core_0.adaptive_ctrl_0.n1705_o[2]\ VPWR VGND _07728_ sg13g2_buf_2
X_14800_ _07727_ _07728_ VPWR VGND _07729_ sg13g2_nor2_1
X_14801_ _07712_ _07723_ _07726_ _07729_ VPWR VGND 
+ _07730_
+ sg13g2_nand4_1
X_14802_ \atbs_core_0.n1386_q\ _07712_ VPWR VGND _07731_ sg13g2_or2_1
X_14803_ \atbs_core_0.comp_upper_sync\ _07718_ _07730_ _07731_ VPWR VGND 
+ _07732_
+ sg13g2_and4_1
X_14804_ _07732_ VPWR VGND _07733_ sg13g2_buf_8
X_14805_ \atbs_core_0.adaptive_mode_uart\ _07653_ VPWR VGND _07734_ sg13g2_nand2_1
X_14806_ _07653_ _07710_ VPWR VGND _07735_ sg13g2_nand2b_1
X_14807_ \atbs_core_0.adaptive_ctrl_0.n1710_o[5]\ VPWR VGND _07736_ sg13g2_buf_8
X_14808_ \atbs_core_0.adaptive_ctrl_0.n1710_o[4]\ VPWR VGND _07737_ sg13g2_buf_4
X_14809_ \atbs_core_0.adaptive_ctrl_0.n1710_o[6]\ VPWR VGND _07738_ sg13g2_buf_4
X_14810_ \atbs_core_0.adaptive_ctrl_0.n1786_q[7]\ VPWR VGND _07739_ sg13g2_buf_2
X_14811_ _07736_ _07737_ _07738_ _07739_ VPWR VGND 
+ _07740_
+ sg13g2_nor4_1
X_14812_ \atbs_core_0.adaptive_ctrl_0.n1710_o[1]\ VPWR VGND _07741_ sg13g2_buf_4
X_14813_ \atbs_core_0.adaptive_ctrl_0.n1710_o[0]\ VPWR VGND _07742_ sg13g2_buf_4
X_14814_ \atbs_core_0.adaptive_ctrl_0.n1710_o[3]\ VPWR VGND _07743_ sg13g2_buf_4
X_14815_ \atbs_core_0.adaptive_ctrl_0.n1710_o[2]\ VPWR VGND _07744_ sg13g2_buf_4
X_14816_ _07741_ _07742_ _07743_ _07744_ VPWR VGND 
+ _07745_
+ sg13g2_nor4_1
X_14817_ _07716_ \atbs_core_0.detection_en\ \atbs_core_0.comp_lower_sync\ VPWR VGND _07746_ sg13g2_nand3b_1
X_14818_ _07734_ _07735_ _07740_ _07745_ _07746_ VPWR 
+ VGND
+ _07747_ sg13g2_a221oi_1
X_14819_ \atbs_core_0.n1387_q\ \atbs_core_0.comp_lower_sync\ VPWR VGND _07748_ sg13g2_nand2_1
X_14820_ _07716_ _07717_ _07712_ _07748_ VPWR VGND 
+ _07749_
+ sg13g2_nor4_1
X_14821_ _00053_ _07747_ _07749_ VPWR VGND _07750_ sg13g2_nor3_2
X_14822_ _07750_ VPWR VGND _07751_ sg13g2_buf_8
X_14823_ _07733_ _07751_ VPWR VGND _07752_ sg13g2_nor2_2
X_14824_ _07752_ VPWR VGND _07753_ sg13g2_buf_8
X_14825_ _07753_ VPWR VGND _07754_ sg13g2_inv_8
X_14826_ _07754_ VPWR VGND _07755_ sg13g2_buf_16
X_14827_ \atbs_core_0.adaptive_ctrl_0.delta_steps[1]\ VPWR VGND _07756_ sg13g2_buf_4
X_14828_ _07756_ VPWR VGND _07757_ sg13g2_inv_1
X_14829_ \atbs_core_0.adaptive_ctrl_0.delta_steps[0]\ VPWR VGND _07758_ sg13g2_buf_1
X_14830_ _07742_ _07758_ VPWR VGND _07759_ sg13g2_nand2b_1
X_14831_ _07741_ _07757_ _07759_ VPWR VGND _07760_ sg13g2_a21oi_1
X_14832_ \atbs_core_0.adaptive_ctrl_0.delta_steps[2]\ VPWR VGND _07761_ sg13g2_buf_4
X_14833_ _07744_ _07761_ VPWR VGND _07762_ sg13g2_nand2b_1
X_14834_ _07741_ _07757_ _07762_ VPWR VGND _07763_ sg13g2_o21ai_1
X_14835_ \atbs_core_0.adaptive_ctrl_0.delta_steps[3]\ VPWR VGND _07764_ sg13g2_buf_4
X_14836_ _07764_ VPWR VGND _07765_ sg13g2_inv_2
X_14837_ _07761_ VPWR VGND _07766_ sg13g2_inv_1
X_14838_ _07743_ _07765_ _07766_ _07744_ VPWR VGND 
+ _07767_
+ sg13g2_a22oi_1
X_14839_ _07760_ _07763_ _07767_ VPWR VGND _07768_ sg13g2_o21ai_1
X_14840_ \atbs_core_0.adaptive_ctrl_0.delta_steps[6]\ VPWR VGND _07769_ sg13g2_buf_4
X_14841_ _07738_ _07769_ VPWR VGND _07770_ sg13g2_nand2b_1
X_14842_ _07769_ _07738_ VPWR VGND _07771_ sg13g2_nand2b_1
X_14843_ \atbs_core_0.adaptive_ctrl_0.delta_steps[4]\ VPWR VGND _07772_ sg13g2_buf_1
X_14844_ _07772_ VPWR VGND _07773_ sg13g2_buf_4
X_14845_ _07737_ _07773_ VPWR VGND _07774_ sg13g2_xnor2_1
X_14846_ _07743_ VPWR VGND _07775_ sg13g2_inv_1
X_14847_ _07736_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ VPWR VGND _07776_ sg13g2_or2_1
X_14848_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ VPWR VGND _07777_ sg13g2_buf_4
X_14849_ _07736_ _07777_ VPWR VGND _07778_ sg13g2_nand2_1
X_14850_ _07775_ _07764_ _07776_ _07778_ _07739_ VPWR 
+ VGND
+ _07779_ sg13g2_a221oi_1
X_14851_ _07770_ _07771_ _07774_ _07779_ VPWR VGND 
+ _07780_
+ sg13g2_and4_1
X_14852_ _07737_ VPWR VGND _07781_ sg13g2_inv_1
X_14853_ _07781_ _07773_ _07777_ VPWR VGND _07782_ sg13g2_o21ai_1
X_14854_ _07781_ _07777_ _07773_ VPWR VGND _07783_ sg13g2_nor3_1
X_14855_ _07736_ _07782_ _07783_ VPWR VGND _07784_ sg13g2_a21o_1
X_14856_ _07739_ _07771_ VPWR VGND _07785_ sg13g2_nand2b_1
X_14857_ _07768_ _07780_ _07784_ _07770_ _07785_ VPWR 
+ VGND
+ _07786_ sg13g2_a221oi_1
X_14858_ _07786_ VPWR VGND _07787_ sg13g2_buf_2
X_14859_ _07787_ VPWR VGND _07788_ sg13g2_buf_4
X_14860_ _07788_ VPWR VGND _07789_ sg13g2_buf_8
X_14861_ _00054_ VPWR VGND _07790_ sg13g2_buf_1
X_14862_ _00052_ _07790_ VPWR VGND _07791_ sg13g2_or2_1
X_14863_ _07715_ _07755_ _07789_ _07791_ VPWR VGND 
+ _07792_
+ sg13g2_nor4_1
X_14864_ _07714_ _07792_ VPWR VGND _07793_ sg13g2_nor2_1
X_14865_ _07793_ VPWR VGND _07794_ sg13g2_buf_1
X_14866_ \atbs_core_0.comp_upper_sync\ _07718_ _07730_ _07731_ VPWR VGND 
+ _07795_
+ sg13g2_nand4_1
X_14867_ _07712_ _07740_ _07745_ VPWR VGND _07796_ sg13g2_nand3_1
X_14868_ \atbs_core_0.n1387_q\ _07712_ _07796_ VPWR VGND _07797_ sg13g2_o21ai_1
X_14869_ _07797_ _07746_ VPWR VGND _07798_ sg13g2_or2_1
X_14870_ _07798_ VPWR VGND _07799_ sg13g2_buf_1
X_14871_ _07795_ _07799_ VPWR VGND _07800_ sg13g2_and2_1
X_14872_ _07800_ VPWR VGND _07801_ sg13g2_buf_1
X_14873_ _07713_ _07801_ VPWR VGND _07802_ sg13g2_nor2_1
X_14874_ _07713_ _07794_ _07802_ VPWR VGND _07803_ sg13g2_a21oi_1
X_14875_ _07709_ _07803_ VPWR VGND _07804_ sg13g2_nor2b_1
X_14876_ _07804_ VPWR VGND _07805_ sg13g2_buf_2
X_14877_ _07805_ VPWR VGND \atbs_core_0.dac_control_0.sync_chain_0.async_i\ sg13g2_inv_1
X_14878_ _07678_ \atbs_core_0.dac_control_0.sync_chain_0.async_i\ VPWR VGND _07806_ sg13g2_nor2_1
X_14879_ _07679_ _07680_ _07806_ VPWR VGND \atbs_core_0.dac_control_0.n1836_o\ sg13g2_a21oi_1
X_14880_ _07713_ VPWR VGND _07807_ sg13g2_buf_1
X_14881_ _07715_ VPWR VGND _07808_ sg13g2_inv_1
X_14882_ _07808_ VPWR VGND _07809_ sg13g2_buf_4
X_14883_ _07728_ VPWR VGND _07810_ sg13g2_inv_1
X_14884_ _07810_ _07761_ VPWR VGND _07811_ sg13g2_nand2_1
X_14885_ _07724_ VPWR VGND _07812_ sg13g2_inv_1
X_14886_ _07725_ _07758_ VPWR VGND _07813_ sg13g2_nor2b_1
X_14887_ _07812_ _07756_ _07813_ VPWR VGND _07814_ sg13g2_o21ai_1
X_14888_ _07812_ _07756_ VPWR VGND _07815_ sg13g2_nand2_1
X_14889_ _07811_ _07814_ _07815_ VPWR VGND _07816_ sg13g2_and3_1
X_14890_ _07777_ _07719_ VPWR VGND _07817_ sg13g2_nor2b_1
X_14891_ _07772_ _07720_ VPWR VGND _07818_ sg13g2_nor2b_1
X_14892_ _07817_ _07818_ VPWR VGND _07819_ sg13g2_nor2_1
X_14893_ _07727_ _07765_ _07766_ _07728_ VPWR VGND 
+ _07820_
+ sg13g2_a22oi_1
X_14894_ _07769_ _07721_ VPWR VGND _07821_ sg13g2_nor2b_1
X_14895_ _07722_ _07821_ VPWR VGND _07822_ sg13g2_nor2_1
X_14896_ _07819_ _07820_ _07822_ VPWR VGND _07823_ sg13g2_nand3_1
X_14897_ _07719_ _07777_ VPWR VGND _07824_ sg13g2_nand2b_1
X_14898_ _07721_ _07769_ VPWR VGND _07825_ sg13g2_nand2b_1
X_14899_ _00055_ _07824_ _07825_ VPWR VGND _07826_ sg13g2_nand3_1
X_14900_ _07722_ _07817_ _07818_ _07821_ VPWR VGND 
+ _07827_
+ sg13g2_nor4_1
X_14901_ _07727_ _07764_ VPWR VGND _07828_ sg13g2_nor2b_1
X_14902_ _07720_ _07773_ VPWR VGND _07829_ sg13g2_nor2b_1
X_14903_ _07817_ _07818_ _07828_ _07829_ VPWR VGND 
+ _07830_
+ sg13g2_or4_1
X_14904_ _07826_ _07822_ _07827_ _07830_ VPWR VGND 
+ _07831_
+ sg13g2_a22oi_1
X_14905_ _07816_ _07823_ _07831_ VPWR VGND _07832_ sg13g2_o21ai_1
X_14906_ _07832_ VPWR VGND _07833_ sg13g2_buf_4
X_14907_ _07833_ VPWR VGND _07834_ sg13g2_buf_8
X_14908_ _07809_ _07834_ VPWR VGND _07835_ sg13g2_nand2_1
X_14909_ _00051_ VPWR VGND _07836_ sg13g2_buf_1
X_14910_ _07733_ _07751_ _07836_ VPWR VGND _07837_ sg13g2_o21ai_1
X_14911_ _07837_ VPWR VGND _07838_ sg13g2_buf_1
X_14912_ _07791_ _07838_ VPWR VGND _07839_ sg13g2_nor2_1
X_14913_ _07835_ _07839_ _07714_ VPWR VGND _07840_ sg13g2_a21oi_1
X_14914_ _07807_ _07840_ _07802_ VPWR VGND _07841_ sg13g2_a21o_1
X_14915_ _07709_ _07841_ VPWR VGND _07842_ sg13g2_nor2_1
X_14916_ _07842_ VPWR VGND _07843_ sg13g2_buf_1
X_14917_ _07843_ VPWR VGND \atbs_core_0.dac_control_1.sync_chain_0.async_i\ sg13g2_inv_1
X_14918_ _07657_ VPWR VGND _07844_ sg13g2_buf_1
X_14919_ \atbs_core_0.dac_control_1.sync_chain_0.async_i\ _07844_ \atbs_core_0.dac_control_1.n1981_o\ VPWR VGND \atbs_core_0.dac_control_1.n1984_o\ sg13g2_mux2_1
X_14920_ _07647_ VPWR VGND _07845_ sg13g2_inv_1
X_14921_ _07645_ VPWR VGND _07846_ sg13g2_inv_1
X_14922_ _07643_ _07644_ VPWR VGND _07847_ sg13g2_nand2_1
X_14923_ _07845_ _07846_ _07847_ VPWR VGND _07848_ sg13g2_nor3_1
X_14924_ _07649_ _07848_ _07637_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3331_o[2]\ sg13g2_mux2_1
X_14925_ \atbs_core_0.atbs_win_length_uart\ VPWR VGND _07849_ sg13g2_buf_1
X_14926_ \atbs_core_0.atbs_max_delta_steps_uart\ _07849_ VPWR VGND _07850_ sg13g2_nor2_1
X_14927_ \atbs_core_0.n1405_q\ VPWR VGND _07851_ sg13g2_buf_1
X_14928_ \atbs_core_0.baudrate_uart\ VPWR VGND _07852_ sg13g2_buf_1
X_14929_ _07851_ _07852_ VPWR VGND _07853_ sg13g2_nor2_1
X_14930_ _07850_ _07853_ VPWR VGND _07854_ sg13g2_and2_1
X_14931_ _07854_ VPWR VGND _07855_ sg13g2_buf_1
X_14932_ \atbs_core_0.n1397_q\ VPWR VGND _07856_ sg13g2_buf_1
X_14933_ \atbs_core_0.n1395_q\ VPWR VGND _07857_ sg13g2_buf_1
X_14934_ \atbs_core_0.n1393_q\ VPWR VGND _07858_ sg13g2_buf_1
X_14935_ \atbs_core_0.analog_trigger_uart\ VPWR VGND _07859_ sg13g2_buf_1
X_14936_ \atbs_core_0.uart_0.rx_data_strb_o\ VPWR VGND _07860_ sg13g2_buf_1
X_14937_ _07859_ _07860_ VPWR VGND _07861_ sg13g2_nand2b_1
X_14938_ _07857_ _07858_ _07861_ VPWR VGND _07862_ sg13g2_nor3_1
X_14939_ _07856_ _07862_ VPWR VGND _07863_ sg13g2_nor2b_1
X_14940_ _07863_ VPWR VGND _07864_ sg13g2_buf_1
X_14941_ \atbs_core_0.n1401_q\ VPWR VGND _07865_ sg13g2_buf_1
X_14942_ \atbs_core_0.n1399_q\ VPWR VGND _07866_ sg13g2_buf_1
X_14943_ _07865_ _07866_ VPWR VGND _07867_ sg13g2_nor2_1
X_14944_ _07864_ _07867_ VPWR VGND _07868_ sg13g2_and2_1
X_14945_ _07855_ _07868_ VPWR VGND _07869_ sg13g2_and2_1
X_14946_ _07869_ VPWR VGND _07870_ sg13g2_buf_1
X_14947_ \atbs_core_0.uart_0.uart_rx_0.n3482_o\ VPWR VGND _07871_ sg13g2_buf_1
X_14948_ \atbs_core_0.uart_0.uart_rx_0.n3480_o\ VPWR VGND _07872_ sg13g2_buf_1
X_14949_ _07872_ VPWR VGND _07873_ sg13g2_inv_1
X_14950_ \atbs_core_0.uart_0.uart_rx_0.n3486_o\ \atbs_core_0.uart_0.uart_rx_0.n3484_o\ VPWR VGND _07874_ sg13g2_nand2b_1
X_14951_ _07874_ VPWR VGND _07875_ sg13g2_buf_1
X_14952_ _07871_ _07873_ _07875_ VPWR VGND _07876_ sg13g2_nor3_1
X_14953_ _07876_ VPWR VGND _07877_ sg13g2_buf_1
X_14954_ \atbs_core_0.uart_0.uart_rx_0.n3472_o\ VPWR VGND _07878_ sg13g2_buf_1
X_14955_ \atbs_core_0.uart_0.uart_rx_0.n3474_o\ VPWR VGND _07879_ sg13g2_buf_1
X_14956_ _07879_ VPWR VGND _07880_ sg13g2_buf_1
X_14957_ \atbs_core_0.uart_0.uart_rx_0.n3476_o\ VPWR VGND _07881_ sg13g2_buf_1
X_14958_ \atbs_core_0.uart_0.uart_rx_0.n3478_o\ VPWR VGND _07882_ sg13g2_buf_1
X_14959_ _07881_ _07882_ VPWR VGND _07883_ sg13g2_nor2_1
X_14960_ _07883_ VPWR VGND _07884_ sg13g2_buf_1
X_14961_ _07880_ _07884_ VPWR VGND _07885_ sg13g2_nand2_1
X_14962_ _07878_ _07885_ VPWR VGND _07886_ sg13g2_nor2_1
X_14963_ _07870_ _07877_ _07886_ VPWR VGND _07887_ sg13g2_nand3_1
X_14964_ \atbs_core_0.n66_o\ _07887_ VPWR VGND _00186_ sg13g2_and2_1
X_14965_ \atbs_core_0.debouncer_0.debounced\ \atbs_core_0.n1383_q\ VPWR VGND _07888_ sg13g2_xor2_1
X_14966_ \atbs_core_0.n1382_q\ \atbs_core_0.debouncer_5.debounced\ VPWR VGND _07889_ sg13g2_xor2_1
X_14967_ \atbs_core_0.n1381_q\ \atbs_core_0.debouncer_3.debounced\ VPWR VGND _07890_ sg13g2_xnor2_1
X_14968_ _07653_ \atbs_core_0.control_mode_d\ VPWR VGND _07891_ sg13g2_xnor2_1
X_14969_ _07710_ \atbs_core_0.adaptive_mode_d\ VPWR VGND _07892_ sg13g2_xnor2_1
X_14970_ _07890_ _07891_ _07892_ VPWR VGND _07893_ sg13g2_nand3_1
X_14971_ _00065_ _07850_ _07877_ VPWR VGND _07894_ sg13g2_nand3_1
X_14972_ _07878_ VPWR VGND _07895_ sg13g2_inv_1
X_14973_ _07895_ _07880_ VPWR VGND _07896_ sg13g2_nor2_1
X_14974_ _07882_ _07881_ VPWR VGND _07897_ sg13g2_nor2b_1
X_14975_ _07897_ VPWR VGND _07898_ sg13g2_buf_1
X_14976_ _07894_ _07896_ _07898_ VPWR VGND _07899_ sg13g2_nand3b_1
X_14977_ _07864_ _07867_ VPWR VGND _07900_ sg13g2_nand2_1
X_14978_ _00064_ _07899_ _07900_ VPWR VGND _07901_ sg13g2_a21oi_1
X_14979_ _07888_ _07889_ _07893_ _07901_ VPWR VGND 
+ _07902_
+ sg13g2_nor4_1
X_14980_ \atbs_core_0.n1412_q[0]\ VPWR VGND _07903_ sg13g2_buf_1
X_14981_ _07685_ _07903_ VPWR VGND _07904_ sg13g2_nand2b_1
X_14982_ _07904_ VPWR VGND _07905_ sg13g2_buf_1
X_14983_ _07681_ _07686_ _07905_ VPWR VGND _07906_ sg13g2_and3_1
X_14984_ _07902_ _07906_ VPWR VGND _07907_ sg13g2_nand2b_1
X_14985_ _00186_ _07907_ VPWR VGND _00185_ sg13g2_and2_1
X_14986_ \atbs_core_0.debouncer_0.debounced\ \atbs_core_0.n1416_q\ _07653_ VPWR VGND _07908_ sg13g2_mux2_1
X_14987_ _07685_ VPWR VGND _07909_ sg13g2_buf_1
X_14988_ _07878_ _07879_ _07884_ VPWR VGND _07910_ sg13g2_nand3_1
X_14989_ _07871_ _07873_ _07875_ _07910_ VPWR VGND 
+ _07911_
+ sg13g2_nor4_1
X_14990_ \atbs_core_0.n72_o\ VPWR VGND _07912_ sg13g2_inv_1
X_14991_ _07912_ \atbs_core_0.n1384_q\ _07908_ VPWR VGND _07913_ sg13g2_o21ai_1
X_14992_ _07870_ _07911_ _07913_ VPWR VGND _07914_ sg13g2_a21oi_1
X_14993_ _07903_ _07681_ VPWR VGND _07915_ sg13g2_nand2b_1
X_14994_ _07914_ _07915_ VPWR VGND _07916_ sg13g2_nor2_1
X_14995_ _07916_ VPWR VGND _07917_ sg13g2_buf_1
X_14996_ _07909_ _07917_ VPWR VGND _07918_ sg13g2_and2_1
X_14997_ _07918_ VPWR VGND _07919_ sg13g2_buf_1
X_14998_ _07908_ _07919_ VPWR VGND _07920_ sg13g2_nand2_1
X_14999_ _00185_ _07920_ VPWR VGND _00188_ sg13g2_and2_1
X_15000_ \atbs_core_0.adaptive_ctrl_0.n1645_o\ VPWR VGND _07921_ sg13g2_buf_1
X_15001_ _07758_ VPWR VGND _07922_ sg13g2_buf_2
X_15002_ _07769_ _07777_ VPWR VGND _07923_ sg13g2_nor2_1
X_15003_ _07773_ _07764_ _07761_ _07756_ VPWR VGND 
+ _07924_
+ sg13g2_nor4_1
X_15004_ _07923_ _07924_ VPWR VGND _07925_ sg13g2_and2_1
X_15005_ _07922_ _07925_ VPWR VGND _07926_ sg13g2_nand2_1
X_15006_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _07921_ _07926_ VPWR VGND _07927_ sg13g2_nand3_1
X_15007_ _07927_ VPWR VGND _07928_ sg13g2_buf_1
X_15008_ _07809_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ _07928_ VPWR VGND _00191_ sg13g2_o21ai_1
X_15009_ _00100_ VPWR VGND _07929_ sg13g2_buf_1
X_15010_ _07929_ VPWR VGND _07930_ sg13g2_buf_1
X_15011_ _07801_ VPWR VGND _07931_ sg13g2_buf_1
X_15012_ _07931_ VPWR VGND _07932_ sg13g2_buf_1
X_15013_ _07930_ _07932_ VPWR VGND _07933_ sg13g2_nand2_1
X_15014_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _07921_ _07933_ VPWR VGND _00192_ sg13g2_mux2_1
X_15015_ \atbs_core_0.adaptive_ctrl_0.n1784_q[0]\ VPWR VGND _07934_ sg13g2_buf_1
X_15016_ _07755_ _07833_ VPWR VGND _07935_ sg13g2_nand2_2
X_15017_ _07753_ VPWR VGND _07936_ sg13g2_buf_4
X_15018_ \atbs_core_0.adaptive_ctrl_0.adaptive_strb\ _07936_ _07789_ VPWR VGND _07937_ sg13g2_nand3_1
X_15019_ _07790_ _07935_ _07937_ VPWR VGND _07938_ sg13g2_o21ai_1
X_15020_ _07836_ _07938_ VPWR VGND _07939_ sg13g2_and2_1
X_15021_ _07939_ VPWR VGND _07940_ sg13g2_buf_1
X_15022_ _07934_ _07940_ VPWR VGND _07941_ sg13g2_nor2b_1
X_15023_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[2]\ VPWR VGND _07942_ sg13g2_a21o_1
X_15024_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ VPWR VGND _07943_ sg13g2_inv_1
X_15025_ _07756_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[1]\ VPWR VGND _07944_ sg13g2_nor2b_1
X_15026_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _07944_ VPWR VGND _07945_ sg13g2_nor2_1
X_15027_ _07761_ _07945_ VPWR VGND _07946_ sg13g2_nor2_1
X_15028_ _07765_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _07944_ _07946_ VPWR 
+ VGND
+ _07947_ sg13g2_a221oi_1
X_15029_ _07764_ _07943_ _07947_ VPWR VGND _07948_ sg13g2_a21oi_1
X_15030_ _07773_ VPWR VGND _07949_ sg13g2_inv_1
X_15031_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _07948_ _07949_ VPWR VGND _07950_ sg13g2_o21ai_1
X_15032_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _07948_ VPWR VGND _07951_ sg13g2_nand2_1
X_15033_ _07950_ _07951_ VPWR VGND _07952_ sg13g2_nand2_1
X_15034_ _07923_ _07942_ _07952_ VPWR VGND _07953_ sg13g2_nand3_1
X_15035_ _07953_ VPWR VGND _07954_ sg13g2_buf_1
X_15036_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[2]\ _07925_ VPWR VGND _07955_ sg13g2_or3_1
X_15037_ \atbs_core_0.adaptive_ctrl_0.n1689_o\ VPWR VGND _07956_ sg13g2_buf_1
X_15038_ _07956_ VPWR VGND _07957_ sg13g2_inv_1
X_15039_ _07954_ _07955_ _07957_ VPWR VGND _07958_ sg13g2_a21oi_1
X_15040_ _07958_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1682_o\ sg13g2_buf_1
X_15041_ _00080_ VPWR VGND _07959_ sg13g2_buf_1
X_15042_ _07959_ _07954_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07960_ sg13g2_nand3b_1
X_15043_ _00151_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ _07960_ VPWR VGND _07961_ sg13g2_o21ai_1
X_15044_ _07919_ _07940_ _07961_ VPWR VGND _07962_ sg13g2_nor3_1
X_15045_ _07941_ _07962_ VPWR VGND _00193_ sg13g2_or2_1
X_15046_ _00084_ _07954_ VPWR VGND _07963_ sg13g2_nand2_1
X_15047_ _07922_ _07954_ _07963_ VPWR VGND _07964_ sg13g2_o21ai_1
X_15048_ _07757_ _07964_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07965_ sg13g2_mux2_1
X_15049_ _07919_ _07940_ VPWR VGND _07966_ sg13g2_or2_1
X_15050_ _07966_ VPWR VGND _07967_ sg13g2_buf_1
X_15051_ \atbs_core_0.adaptive_ctrl_0.n1784_q[1]\ VPWR VGND _07968_ sg13g2_buf_1
X_15052_ _07968_ _07940_ VPWR VGND _07969_ sg13g2_nand2_1
X_15053_ _07965_ _07967_ _07969_ VPWR VGND _00194_ sg13g2_o21ai_1
X_15054_ _07959_ _00082_ _07954_ VPWR VGND _07970_ sg13g2_mux2_1
X_15055_ _07766_ _07970_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07971_ sg13g2_mux2_1
X_15056_ \atbs_core_0.adaptive_ctrl_0.n1784_q[2]\ VPWR VGND _07972_ sg13g2_buf_1
X_15057_ _07972_ _07940_ VPWR VGND _07973_ sg13g2_nand2_1
X_15058_ _07967_ _07971_ _07973_ VPWR VGND _00195_ sg13g2_o21ai_1
X_15059_ _00084_ _00088_ _07954_ VPWR VGND _07974_ sg13g2_mux2_1
X_15060_ _07765_ _07974_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07975_ sg13g2_mux2_1
X_15061_ \atbs_core_0.adaptive_ctrl_0.n1784_q[3]\ VPWR VGND _07976_ sg13g2_buf_1
X_15062_ _07976_ _07940_ VPWR VGND _07977_ sg13g2_nand2_1
X_15063_ _07967_ _07975_ _07977_ VPWR VGND _00196_ sg13g2_o21ai_1
X_15064_ _00082_ _00086_ _07954_ VPWR VGND _07978_ sg13g2_mux2_1
X_15065_ _07949_ _07978_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07979_ sg13g2_mux2_1
X_15066_ \atbs_core_0.adaptive_ctrl_0.n1784_q[4]\ VPWR VGND _07980_ sg13g2_buf_1
X_15067_ _07980_ _07940_ VPWR VGND _07981_ sg13g2_nand2_1
X_15068_ _07967_ _07979_ _07981_ VPWR VGND _00197_ sg13g2_o21ai_1
X_15069_ _07777_ VPWR VGND _07982_ sg13g2_inv_1
X_15070_ _00088_ _00090_ _07954_ VPWR VGND _07983_ sg13g2_mux2_1
X_15071_ _07982_ _07983_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07984_ sg13g2_mux2_1
X_15072_ \atbs_core_0.adaptive_ctrl_0.n1784_q[5]\ VPWR VGND _07985_ sg13g2_buf_1
X_15073_ _07985_ _07940_ VPWR VGND _07986_ sg13g2_nand2_1
X_15074_ _07967_ _07984_ _07986_ VPWR VGND _00198_ sg13g2_o21ai_1
X_15075_ \atbs_core_0.adaptive_ctrl_0.n1682_o\ VPWR VGND _07987_ sg13g2_inv_1
X_15076_ _00086_ _07957_ _07954_ VPWR VGND _07988_ sg13g2_nor3_1
X_15077_ _07769_ _07987_ _07988_ VPWR VGND _07989_ sg13g2_a21oi_1
X_15078_ \atbs_core_0.adaptive_ctrl_0.n1784_q[6]\ _07940_ VPWR VGND _07990_ sg13g2_nand2_1
X_15079_ _07967_ _07989_ _07990_ VPWR VGND _00199_ sg13g2_o21ai_1
X_15080_ _07909_ _07917_ VPWR VGND _07991_ sg13g2_nand2_1
X_15081_ _07991_ VPWR VGND _07992_ sg13g2_buf_1
X_15082_ _07922_ _07956_ VPWR VGND _07993_ sg13g2_nand2_1
X_15083_ _07956_ _00152_ _07993_ VPWR VGND _07994_ sg13g2_o21ai_1
X_15084_ _07992_ _07994_ VPWR VGND _00200_ sg13g2_nand2_1
X_15085_ _07919_ VPWR VGND _07995_ sg13g2_buf_1
X_15086_ _07957_ VPWR VGND _07996_ sg13g2_buf_1
X_15087_ _07757_ _07996_ VPWR VGND _07997_ sg13g2_nor2_1
X_15088_ _07968_ _07996_ _07997_ VPWR VGND _07998_ sg13g2_a21oi_1
X_15089_ _07995_ _07998_ VPWR VGND _00201_ sg13g2_nor2_1
X_15090_ _07766_ _07996_ VPWR VGND _07999_ sg13g2_nor2_1
X_15091_ _07972_ _07996_ _07999_ VPWR VGND _08000_ sg13g2_a21oi_1
X_15092_ _07995_ _08000_ VPWR VGND _00202_ sg13g2_nor2_1
X_15093_ _07765_ _07996_ VPWR VGND _08001_ sg13g2_nor2_1
X_15094_ _07976_ _07996_ _08001_ VPWR VGND _08002_ sg13g2_a21oi_1
X_15095_ _07995_ _08002_ VPWR VGND _00203_ sg13g2_nor2_1
X_15096_ _07949_ _07957_ VPWR VGND _08003_ sg13g2_nor2_1
X_15097_ _07980_ _07996_ _08003_ VPWR VGND _08004_ sg13g2_a21oi_1
X_15098_ _07995_ _08004_ VPWR VGND _00204_ sg13g2_nor2_1
X_15099_ _07982_ _07957_ VPWR VGND _08005_ sg13g2_nor2_1
X_15100_ _07985_ _07996_ _08005_ VPWR VGND _08006_ sg13g2_a21oi_1
X_15101_ _07995_ _08006_ VPWR VGND _00205_ sg13g2_nor2_1
X_15102_ _07769_ _07956_ VPWR VGND _08007_ sg13g2_and2_1
X_15103_ \atbs_core_0.adaptive_ctrl_0.n1784_q[6]\ _07996_ _08007_ VPWR VGND _08008_ sg13g2_a21oi_1
X_15104_ _07995_ _08008_ VPWR VGND _00206_ sg13g2_nor2_1
X_15105_ _07909_ VPWR VGND _08009_ sg13g2_buf_1
X_15106_ _07715_ _07733_ _07751_ VPWR VGND _08010_ sg13g2_nor3_1
X_15107_ _08010_ VPWR VGND _08011_ sg13g2_buf_4
X_15108_ _07742_ _07788_ _08011_ VPWR VGND _08012_ sg13g2_and3_1
X_15109_ _08012_ VPWR VGND _08013_ sg13g2_buf_2
X_15110_ _07725_ _07809_ _07755_ _07833_ VPWR VGND 
+ _08014_
+ sg13g2_and4_1
X_15111_ _08014_ VPWR VGND _08015_ sg13g2_buf_2
X_15112_ _08013_ _08015_ VPWR VGND _08016_ sg13g2_nor2_1
X_15113_ _07809_ _07755_ _07833_ VPWR VGND _08017_ sg13g2_nand3_1
X_15114_ _08017_ VPWR VGND _08018_ sg13g2_buf_8
X_15115_ _07787_ _08011_ VPWR VGND _08019_ sg13g2_nand2_1
X_15116_ _08019_ VPWR VGND _08020_ sg13g2_buf_2
X_15117_ _07790_ _07715_ \atbs_core_0.adaptive_ctrl_0.n1781_q\ VPWR VGND _08021_ sg13g2_or3_1
X_15118_ _08021_ VPWR VGND _08022_ sg13g2_buf_1
X_15119_ _07733_ _07751_ _08022_ VPWR VGND _08023_ sg13g2_nor3_1
X_15120_ _07789_ _08023_ _07934_ VPWR VGND _08024_ sg13g2_nand3b_1
X_15121_ _07922_ _08018_ _08020_ _08024_ VPWR VGND 
+ _08025_
+ sg13g2_nand4_1
X_15122_ _07922_ VPWR VGND _08026_ sg13g2_inv_1
X_15123_ _08024_ _08026_ VPWR VGND _08027_ sg13g2_nand2b_1
X_15124_ _08016_ _08025_ _08027_ VPWR VGND _08028_ sg13g2_nand3_1
X_15125_ _08028_ VPWR VGND _08029_ sg13g2_buf_1
X_15126_ _07725_ _08029_ VPWR VGND _08030_ sg13g2_xor2_1
X_15127_ _07794_ VPWR VGND _08031_ sg13g2_buf_1
X_15128_ _00153_ _08031_ VPWR VGND _08032_ sg13g2_nor2_1
X_15129_ _08009_ _07917_ _08030_ _08031_ _08032_ VPWR 
+ VGND
+ _00207_ sg13g2_a221oi_1
X_15130_ _07792_ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ VPWR VGND _08033_ sg13g2_nand2b_1
X_15131_ _08033_ VPWR VGND _08034_ sg13g2_buf_1
X_15132_ _07724_ _08034_ VPWR VGND _08035_ sg13g2_nand2_1
X_15133_ _00081_ VPWR VGND _08036_ sg13g2_buf_1
X_15134_ _08036_ VPWR VGND _08037_ sg13g2_inv_1
X_15135_ _07753_ _07787_ _07959_ VPWR VGND _08038_ sg13g2_a21oi_1
X_15136_ _07741_ VPWR VGND _08039_ sg13g2_inv_1
X_15137_ _08039_ _07715_ _07733_ _07751_ VPWR VGND 
+ _08040_
+ sg13g2_nor4_1
X_15138_ _07809_ _07959_ VPWR VGND _08041_ sg13g2_nor2_1
X_15139_ _07787_ _08040_ _08041_ VPWR VGND _08042_ sg13g2_a21o_1
X_15140_ _07935_ _08038_ _08042_ VPWR VGND _08043_ sg13g2_a21oi_1
X_15141_ _08043_ VPWR VGND _08044_ sg13g2_buf_4
X_15142_ _07819_ _07820_ _07822_ VPWR VGND _08045_ sg13g2_and3_1
X_15143_ _07811_ _07814_ _07815_ VPWR VGND _08046_ sg13g2_nand3_1
X_15144_ _07830_ _07827_ VPWR VGND _08047_ sg13g2_and2_1
X_15145_ _07826_ _07822_ _08045_ _08046_ _08047_ VPWR 
+ VGND
+ _08048_ sg13g2_a221oi_1
X_15146_ _08048_ VPWR VGND _08049_ sg13g2_buf_2
X_15147_ _07715_ _07753_ _08049_ VPWR VGND _08050_ sg13g2_nor3_2
X_15148_ _08050_ VPWR VGND _08051_ sg13g2_buf_4
X_15149_ _07733_ _07751_ _08022_ VPWR VGND _08052_ sg13g2_or3_1
X_15150_ _08052_ VPWR VGND _08053_ sg13g2_buf_2
X_15151_ _07788_ _08053_ VPWR VGND _08054_ sg13g2_nor2_1
X_15152_ _08054_ VPWR VGND _08055_ sg13g2_buf_4
X_15153_ _08051_ _08055_ VPWR VGND _08056_ sg13g2_nor2_1
X_15154_ _07788_ _08023_ VPWR VGND _08057_ sg13g2_nand2b_1
X_15155_ _08057_ VPWR VGND _08058_ sg13g2_buf_2
X_15156_ _07922_ _07934_ VPWR VGND _08059_ sg13g2_nand2_1
X_15157_ _07756_ _07968_ VPWR VGND _08060_ sg13g2_xor2_1
X_15158_ _08059_ _08060_ VPWR VGND _08061_ sg13g2_xnor2_1
X_15159_ _08058_ _08061_ VPWR VGND _08062_ sg13g2_nor2_1
X_15160_ _08044_ _08056_ _08062_ VPWR VGND _08063_ sg13g2_a21o_1
X_15161_ _07755_ _07789_ VPWR VGND _08064_ sg13g2_nor2_1
X_15162_ _08022_ _08061_ VPWR VGND _08065_ sg13g2_nor2_1
X_15163_ _08064_ _08065_ _08044_ _08058_ _08037_ VPWR 
+ VGND
+ _08066_ sg13g2_a221oi_1
X_15164_ _08037_ _08063_ _08066_ VPWR VGND _08067_ sg13g2_a21oi_1
X_15165_ _07725_ _07838_ VPWR VGND _08068_ sg13g2_xnor2_1
X_15166_ _08029_ _08067_ _08068_ VPWR VGND _08069_ sg13g2_and3_1
X_15167_ _08029_ _08068_ _08067_ VPWR VGND _08070_ sg13g2_a21oi_1
X_15168_ _08069_ _08070_ _08031_ VPWR VGND _08071_ sg13g2_o21ai_1
X_15169_ _08035_ _08071_ _07995_ VPWR VGND _00208_ sg13g2_a21oi_1
X_15170_ _00154_ _08034_ VPWR VGND _08072_ sg13g2_nand2_1
X_15171_ _07755_ VPWR VGND spike_o sg13g2_buf_8
X_15172_ _08037_ _08051_ _08055_ VPWR VGND _08073_ sg13g2_a21oi_1
X_15173_ _07836_ spike_o _08044_ _08073_ _08062_ VPWR 
+ VGND
+ _08074_ sg13g2_a221oi_1
X_15174_ _07959_ _08018_ _08020_ VPWR VGND _08075_ sg13g2_nand3b_1
X_15175_ _08037_ _08051_ VPWR VGND _08076_ sg13g2_nand2_1
X_15176_ _08075_ _08076_ _07725_ VPWR VGND _08077_ sg13g2_a21oi_1
X_15177_ _07836_ spike_o VPWR VGND _08078_ sg13g2_and2_1
X_15178_ _08078_ VPWR VGND _08079_ sg13g2_buf_1
X_15179_ _07725_ _08037_ _08079_ VPWR VGND _08080_ sg13g2_a21oi_1
X_15180_ _07726_ _08074_ _08077_ _08080_ VPWR VGND 
+ _08081_
+ sg13g2_or4_1
X_15181_ _08025_ _08027_ VPWR VGND _08082_ sg13g2_and2_1
X_15182_ _07724_ _08036_ VPWR VGND _08083_ sg13g2_nor2_1
X_15183_ _07726_ _08083_ VPWR VGND _08084_ sg13g2_nor2_1
X_15184_ _08016_ _08082_ _08074_ _08084_ VPWR VGND 
+ _08085_
+ sg13g2_a22oi_1
X_15185_ _08063_ _08083_ _08066_ VPWR VGND _08086_ sg13g2_a21o_1
X_15186_ _07838_ _08029_ VPWR VGND _08087_ sg13g2_nand2_1
X_15187_ _08081_ _08085_ _08086_ _08087_ VPWR VGND 
+ _08088_
+ sg13g2_a22oi_1
X_15188_ _07922_ _08018_ _08020_ VPWR VGND _08089_ sg13g2_nand3_1
X_15189_ _08089_ VPWR VGND _08090_ sg13g2_buf_2
X_15190_ _08037_ _08050_ _08038_ _07935_ _08042_ VPWR 
+ VGND
+ _08091_ sg13g2_a221oi_1
X_15191_ _08091_ VPWR VGND _08092_ sg13g2_buf_4
X_15192_ _08016_ _08090_ _08092_ VPWR VGND _08093_ sg13g2_nand3_1
X_15193_ _08093_ VPWR VGND _08094_ sg13g2_buf_2
X_15194_ _00084_ _08018_ _08020_ VPWR VGND _08095_ sg13g2_nand3b_1
X_15195_ _08095_ VPWR VGND _08096_ sg13g2_buf_4
X_15196_ _07744_ _07789_ _08011_ VPWR VGND _08097_ sg13g2_nand3_1
X_15197_ _07728_ _07809_ _07755_ _07834_ VPWR VGND 
+ _08098_
+ sg13g2_nand4_1
X_15198_ _08097_ _08098_ VPWR VGND _08099_ sg13g2_and2_1
X_15199_ _08099_ VPWR VGND _08100_ sg13g2_buf_1
X_15200_ _08096_ _08100_ _08055_ VPWR VGND _08101_ sg13g2_a21oi_1
X_15201_ _07761_ _07972_ VPWR VGND _08102_ sg13g2_xor2_1
X_15202_ _07756_ _07968_ _07934_ _07922_ VPWR VGND 
+ _08103_
+ sg13g2_a22oi_1
X_15203_ _07756_ _07968_ VPWR VGND _08104_ sg13g2_nor2_1
X_15204_ _08103_ _08104_ VPWR VGND _08105_ sg13g2_nor2_1
X_15205_ _08102_ _08105_ VPWR VGND _08106_ sg13g2_xnor2_1
X_15206_ _08106_ VPWR VGND _08107_ sg13g2_buf_1
X_15207_ _07922_ _07934_ VPWR VGND _08108_ sg13g2_xor2_1
X_15208_ _08061_ _08108_ VPWR VGND _08109_ sg13g2_nor2_1
X_15209_ _08107_ _08109_ VPWR VGND _08110_ sg13g2_nor2_1
X_15210_ _08094_ _08101_ _08110_ _08055_ VPWR VGND 
+ _08111_
+ sg13g2_a22oi_1
X_15211_ _08096_ _08100_ VPWR VGND _08112_ sg13g2_and2_1
X_15212_ _08112_ VPWR VGND _08113_ sg13g2_buf_1
X_15213_ _08058_ _08096_ _08100_ VPWR VGND _08114_ sg13g2_and3_1
X_15214_ _08016_ _08090_ _08092_ VPWR VGND _08115_ sg13g2_and3_1
X_15215_ _08115_ VPWR VGND _08116_ sg13g2_buf_2
X_15216_ _08107_ _08109_ VPWR VGND _08117_ sg13g2_and2_1
X_15217_ _08117_ VPWR VGND _08118_ sg13g2_buf_1
X_15218_ _08055_ _08118_ VPWR VGND _08119_ sg13g2_and2_1
X_15219_ _08079_ _08113_ _08114_ _08116_ _08119_ VPWR 
+ VGND
+ _08120_ sg13g2_a221oi_1
X_15220_ _08079_ _08111_ _08120_ VPWR VGND _08121_ sg13g2_o21ai_1
X_15221_ _07810_ _08121_ VPWR VGND _08122_ sg13g2_xnor2_1
X_15222_ _08088_ _08122_ VPWR VGND _08123_ sg13g2_xnor2_1
X_15223_ _08031_ _08123_ VPWR VGND _08124_ sg13g2_nand2_1
X_15224_ _08072_ _08124_ _07995_ VPWR VGND _00209_ sg13g2_a21oi_1
X_15225_ _08088_ _08121_ VPWR VGND _08125_ sg13g2_and2_1
X_15226_ _08125_ VPWR VGND _08126_ sg13g2_buf_1
X_15227_ _08088_ _08121_ VPWR VGND _08127_ sg13g2_or2_1
X_15228_ _08127_ VPWR VGND _08128_ sg13g2_buf_1
X_15229_ _07728_ _08126_ _08128_ VPWR VGND _08129_ sg13g2_o21ai_1
X_15230_ _08079_ _08119_ VPWR VGND _08130_ sg13g2_or2_1
X_15231_ _08116_ _08114_ _08130_ VPWR VGND _08131_ sg13g2_a21o_1
X_15232_ _00082_ _08018_ _08020_ VPWR VGND _08132_ sg13g2_nand3b_1
X_15233_ _08132_ VPWR VGND _08133_ sg13g2_buf_2
X_15234_ _07743_ _07788_ _08011_ VPWR VGND _08134_ sg13g2_nand3_1
X_15235_ _07727_ _07809_ _07755_ _07833_ VPWR VGND 
+ _08135_
+ sg13g2_nand4_1
X_15236_ _08134_ _08135_ VPWR VGND _08136_ sg13g2_and2_1
X_15237_ _08136_ VPWR VGND _08137_ sg13g2_buf_1
X_15238_ _08133_ _08137_ VPWR VGND _08138_ sg13g2_and2_1
X_15239_ _08138_ VPWR VGND _08139_ sg13g2_buf_1
X_15240_ _07761_ _07972_ VPWR VGND _08140_ sg13g2_nor2_1
X_15241_ _08103_ _08104_ _08140_ VPWR VGND _08141_ sg13g2_nor3_1
X_15242_ _07761_ _07972_ _08141_ VPWR VGND _08142_ sg13g2_a21oi_1
X_15243_ _07764_ _07976_ VPWR VGND _08143_ sg13g2_xor2_1
X_15244_ _08142_ _08143_ VPWR VGND _08144_ sg13g2_xnor2_1
X_15245_ _07789_ _08053_ _08144_ VPWR VGND _08145_ sg13g2_nor3_2
X_15246_ _08058_ _08139_ _08145_ VPWR VGND _08146_ sg13g2_a21o_1
X_15247_ _08131_ _08146_ VPWR VGND _08147_ sg13g2_xor2_1
X_15248_ _07727_ _08147_ VPWR VGND _08148_ sg13g2_xnor2_1
X_15249_ _08129_ _08148_ VPWR VGND _08149_ sg13g2_xnor2_1
X_15250_ _00155_ _08031_ VPWR VGND _08150_ sg13g2_nor2_1
X_15251_ _08009_ _07917_ _08149_ _08031_ _08150_ VPWR 
+ VGND
+ _00210_ sg13g2_a221oi_1
X_15252_ _07727_ VPWR VGND _08151_ sg13g2_inv_1
X_15253_ _08151_ _08147_ VPWR VGND _08152_ sg13g2_nand2_1
X_15254_ _08151_ _08147_ _07810_ VPWR VGND _08153_ sg13g2_a21oi_1
X_15255_ _08151_ _08147_ VPWR VGND _08154_ sg13g2_nor2_1
X_15256_ _08126_ _08152_ _08153_ _08128_ _08154_ VPWR 
+ VGND
+ _08155_ sg13g2_a221oi_1
X_15257_ _08155_ VPWR VGND _08156_ sg13g2_buf_1
X_15258_ _07720_ VPWR VGND _08157_ sg13g2_inv_1
X_15259_ _07773_ _07980_ VPWR VGND _08158_ sg13g2_xnor2_1
X_15260_ _07764_ _07976_ VPWR VGND _08159_ sg13g2_nand2_1
X_15261_ _07764_ _07976_ VPWR VGND _08160_ sg13g2_nor2_1
X_15262_ _08142_ _08159_ _08160_ VPWR VGND _08161_ sg13g2_a21oi_1
X_15263_ _08158_ _08161_ VPWR VGND _08162_ sg13g2_xnor2_1
X_15264_ _07788_ _08011_ VPWR VGND _08163_ sg13g2_and2_1
X_15265_ _08163_ VPWR VGND _08164_ sg13g2_buf_2
X_15266_ _00088_ _08051_ _08164_ VPWR VGND _08165_ sg13g2_nor3_1
X_15267_ _07737_ _07788_ _08011_ VPWR VGND _08166_ sg13g2_nand3_1
X_15268_ _08157_ _08018_ _08166_ VPWR VGND _08167_ sg13g2_o21ai_1
X_15269_ _08167_ VPWR VGND _08168_ sg13g2_buf_1
X_15270_ _08165_ _08168_ VPWR VGND _08169_ sg13g2_or2_1
X_15271_ _08162_ _08169_ _08058_ VPWR VGND _08170_ sg13g2_mux2_1
X_15272_ _08170_ VPWR VGND _08171_ sg13g2_buf_1
X_15273_ _08058_ _08116_ _08113_ _08139_ VPWR VGND 
+ _08172_
+ sg13g2_nand4_1
X_15274_ _08172_ VPWR VGND _08173_ sg13g2_buf_1
X_15275_ _08118_ _08145_ _08079_ VPWR VGND _08174_ sg13g2_a21oi_1
X_15276_ _08173_ _08174_ VPWR VGND _08175_ sg13g2_nand2_1
X_15277_ _08171_ _08175_ VPWR VGND _08176_ sg13g2_xor2_1
X_15278_ _08157_ _08176_ VPWR VGND _08177_ sg13g2_xnor2_1
X_15279_ _08156_ _08177_ VPWR VGND _08178_ sg13g2_xnor2_1
X_15280_ _00156_ _08031_ VPWR VGND _08179_ sg13g2_nor2_1
X_15281_ _08009_ _07917_ _08178_ _08031_ _08179_ VPWR 
+ VGND
+ _00211_ sg13g2_a221oi_1
X_15282_ _08126_ _08152_ _08153_ _08128_ VPWR VGND 
+ _08180_
+ sg13g2_a22oi_1
X_15283_ _08154_ _08180_ VPWR VGND _08181_ sg13g2_nand2b_1
X_15284_ _08176_ VPWR VGND _08182_ sg13g2_inv_1
X_15285_ _08156_ _08182_ _08157_ VPWR VGND _08183_ sg13g2_o21ai_1
X_15286_ _08181_ _08176_ _08183_ VPWR VGND _08184_ sg13g2_o21ai_1
X_15287_ _07719_ VPWR VGND _08185_ sg13g2_inv_1
X_15288_ _07761_ _07972_ _07980_ _07773_ VPWR VGND 
+ _08186_
+ sg13g2_a22oi_1
X_15289_ _07976_ _08186_ VPWR VGND _08187_ sg13g2_nand2b_1
X_15290_ _07765_ _08186_ VPWR VGND _08188_ sg13g2_nand2_1
X_15291_ _08187_ _08188_ _08141_ VPWR VGND _08189_ sg13g2_a21oi_1
X_15292_ _07773_ _07980_ VPWR VGND _08190_ sg13g2_nand2_1
X_15293_ _07773_ _07980_ VPWR VGND _08191_ sg13g2_nor2_1
X_15294_ _08160_ _08190_ _08191_ VPWR VGND _08192_ sg13g2_a21oi_1
X_15295_ _08189_ _08192_ VPWR VGND _08193_ sg13g2_nand2b_1
X_15296_ _07777_ _07985_ VPWR VGND _08194_ sg13g2_xor2_1
X_15297_ _08193_ _08194_ VPWR VGND _08195_ sg13g2_xnor2_1
X_15298_ _08058_ _08195_ VPWR VGND _08196_ sg13g2_or2_1
X_15299_ _08196_ VPWR VGND _08197_ sg13g2_buf_1
X_15300_ _07719_ _08051_ _08164_ _07736_ VPWR VGND 
+ _08198_
+ sg13g2_a22oi_1
X_15301_ _00086_ _08018_ _08020_ VPWR VGND _08199_ sg13g2_nand3b_1
X_15302_ _08058_ _08198_ _08199_ VPWR VGND _08200_ sg13g2_nand3_1
X_15303_ _08200_ VPWR VGND _08201_ sg13g2_buf_2
X_15304_ _08197_ _08201_ VPWR VGND _08202_ sg13g2_nand2_1
X_15305_ _08174_ _08202_ VPWR VGND _08203_ sg13g2_and2_1
X_15306_ _08171_ _08202_ VPWR VGND _08204_ sg13g2_and2_1
X_15307_ _07838_ _08171_ _08173_ _08174_ _08202_ VPWR 
+ VGND
+ _08205_ sg13g2_a221oi_1
X_15308_ _08173_ _08203_ _08204_ _07838_ _08205_ VPWR 
+ VGND
+ _08206_ sg13g2_a221oi_1
X_15309_ _08206_ VPWR VGND _08207_ sg13g2_buf_1
X_15310_ _08185_ _08207_ VPWR VGND _08208_ sg13g2_xnor2_1
X_15311_ _08184_ _08208_ VPWR VGND _08209_ sg13g2_xnor2_1
X_15312_ _00157_ _07794_ _07992_ VPWR VGND _08210_ sg13g2_o21ai_1
X_15313_ _08031_ _08209_ _08210_ VPWR VGND _00212_ sg13g2_a21oi_1
X_15314_ _08173_ _08203_ _08204_ _07838_ VPWR VGND 
+ _08211_
+ sg13g2_a22oi_1
X_15315_ _08205_ _08211_ VPWR VGND _08212_ sg13g2_nand2b_1
X_15316_ _08157_ _08182_ _08212_ _08185_ _08156_ VPWR 
+ VGND
+ _08213_ sg13g2_a221oi_1
X_15317_ _07719_ _08207_ VPWR VGND _08214_ sg13g2_nand2_1
X_15318_ _07720_ _08176_ _08207_ VPWR VGND _08215_ sg13g2_nand3_1
X_15319_ _07719_ _07720_ _08176_ VPWR VGND _08216_ sg13g2_nand3_1
X_15320_ _08214_ _08215_ _08216_ VPWR VGND _08217_ sg13g2_nand3_1
X_15321_ _08213_ _08217_ VPWR VGND _08218_ sg13g2_nor2_1
X_15322_ _00091_ VPWR VGND _08219_ sg13g2_buf_1
X_15323_ _00092_ VPWR VGND _08220_ sg13g2_inv_1
X_15324_ _08220_ _07936_ _07789_ VPWR VGND _08221_ sg13g2_nand3_1
X_15325_ _08219_ _07935_ _08221_ VPWR VGND _08222_ sg13g2_o21ai_1
X_15326_ _00090_ _08051_ _08164_ VPWR VGND _08223_ sg13g2_nor3_1
X_15327_ _07809_ _08222_ _08223_ VPWR VGND _08224_ sg13g2_a21oi_1
X_15328_ _07777_ _07985_ VPWR VGND _08225_ sg13g2_nand2_1
X_15329_ _07777_ _07985_ VPWR VGND _08226_ sg13g2_nor2_1
X_15330_ _08193_ _08225_ _08226_ VPWR VGND _08227_ sg13g2_a21oi_1
X_15331_ _07769_ \atbs_core_0.adaptive_ctrl_0.n1784_q[6]\ VPWR VGND _08228_ sg13g2_xnor2_1
X_15332_ _08227_ _08228_ VPWR VGND _08229_ sg13g2_xnor2_1
X_15333_ _08058_ _08229_ VPWR VGND _08230_ sg13g2_nor2_1
X_15334_ _08058_ _08224_ _08230_ VPWR VGND _08231_ sg13g2_a21o_1
X_15335_ _08231_ VPWR VGND _08232_ sg13g2_buf_1
X_15336_ _08118_ _08145_ VPWR VGND _08233_ sg13g2_nand2_1
X_15337_ _08173_ _08233_ _08197_ _08201_ _08171_ VPWR 
+ VGND
+ _08234_ sg13g2_a221oi_1
X_15338_ _08079_ _08234_ VPWR VGND _08235_ sg13g2_nor2_1
X_15339_ _08232_ _08235_ VPWR VGND _08236_ sg13g2_xnor2_1
X_15340_ _08219_ _08236_ VPWR VGND _08237_ sg13g2_xnor2_1
X_15341_ _08218_ _08237_ VPWR VGND _08238_ sg13g2_xnor2_1
X_15342_ _07721_ _07794_ _07992_ VPWR VGND _08239_ sg13g2_o21ai_1
X_15343_ _08031_ _08238_ _08239_ VPWR VGND _00213_ sg13g2_a21oi_1
X_15344_ _07721_ VPWR VGND _08240_ sg13g2_inv_1
X_15345_ _07721_ _08219_ VPWR VGND _08241_ sg13g2_or2_1
X_15346_ _08232_ _08234_ _08079_ VPWR VGND _08242_ sg13g2_a21oi_1
X_15347_ _00055_ _08242_ VPWR VGND _08243_ sg13g2_xor2_1
X_15348_ _08240_ _08241_ _08243_ VPWR VGND _08244_ sg13g2_mux2_1
X_15349_ _08219_ _08236_ _08243_ VPWR VGND _08245_ sg13g2_nand3_1
X_15350_ _08236_ _08244_ _08245_ VPWR VGND _08246_ sg13g2_o21ai_1
X_15351_ _07722_ _08034_ VPWR VGND _08247_ sg13g2_nand2b_1
X_15352_ _08034_ _08246_ _08247_ VPWR VGND _08248_ sg13g2_o21ai_1
X_15353_ _08034_ _07919_ _08237_ _08243_ VPWR VGND 
+ _08249_
+ sg13g2_or4_1
X_15354_ _08240_ _08236_ _07794_ VPWR VGND _08250_ sg13g2_o21ai_1
X_15355_ _08250_ _08243_ _07992_ VPWR VGND _08251_ sg13g2_nand3b_1
X_15356_ _08249_ _08251_ _08218_ VPWR VGND _08252_ sg13g2_mux2_1
X_15357_ _07919_ _08248_ _08252_ VPWR VGND _00214_ sg13g2_o21ai_1
X_15358_ _07790_ _07715_ \atbs_core_0.adaptive_ctrl_0.n1781_q\ VPWR VGND _08253_ sg13g2_nor3_1
X_15359_ _07934_ _08253_ VPWR VGND _08254_ sg13g2_nand2_1
X_15360_ _07753_ _07834_ _08254_ VPWR VGND _08255_ sg13g2_nor3_1
X_15361_ _08026_ _08051_ _08164_ _08255_ VPWR VGND 
+ _08256_
+ sg13g2_or4_1
X_15362_ _07922_ _07753_ _07834_ _08254_ VPWR VGND 
+ _08257_
+ sg13g2_nor4_1
X_15363_ _08013_ _08015_ _08257_ VPWR VGND _08258_ sg13g2_nor3_1
X_15364_ _08256_ _08258_ VPWR VGND _08259_ sg13g2_and2_1
X_15365_ _08259_ VPWR VGND _08260_ sg13g2_buf_1
X_15366_ _07742_ _08260_ VPWR VGND _08261_ sg13g2_xnor2_1
X_15367_ _07840_ VPWR VGND _08262_ sg13g2_buf_1
X_15368_ _00158_ _08262_ VPWR VGND _08263_ sg13g2_nor2_1
X_15369_ _08009_ _07917_ _08261_ _08262_ _08263_ VPWR 
+ VGND
+ _00215_ sg13g2_a221oi_1
X_15370_ _08011_ VPWR VGND _08264_ sg13g2_buf_1
X_15371_ _07742_ _08264_ VPWR VGND _08265_ sg13g2_xnor2_1
X_15372_ _08260_ _08265_ VPWR VGND _08266_ sg13g2_nor2_1
X_15373_ _07936_ _07834_ VPWR VGND _08267_ sg13g2_nor2_1
X_15374_ _07715_ _08036_ VPWR VGND _08268_ sg13g2_nor2_1
X_15375_ _08253_ _08268_ _07834_ VPWR VGND _08269_ sg13g2_mux2_1
X_15376_ spike_o _08269_ VPWR VGND _08270_ sg13g2_nand2_1
X_15377_ _08065_ _08267_ _08270_ _08044_ VPWR VGND 
+ _08271_
+ sg13g2_a22oi_1
X_15378_ _07741_ _08271_ VPWR VGND _08272_ sg13g2_xnor2_1
X_15379_ _08266_ _08272_ VPWR VGND _08273_ sg13g2_xnor2_1
X_15380_ _00159_ _08262_ VPWR VGND _08274_ sg13g2_nor2_1
X_15381_ _08009_ _07917_ _08273_ _08262_ _08274_ VPWR 
+ VGND
+ _00216_ sg13g2_a221oi_1
X_15382_ _07835_ _07839_ _07714_ VPWR VGND _08275_ sg13g2_a21o_1
X_15383_ _08275_ VPWR VGND _08276_ sg13g2_buf_1
X_15384_ _07809_ _07753_ VPWR VGND _08277_ sg13g2_nand2_1
X_15385_ _08277_ VPWR VGND _08278_ sg13g2_buf_1
X_15386_ _08026_ _07789_ _08278_ VPWR VGND _08279_ sg13g2_nor3_1
X_15387_ _08039_ _08013_ _08279_ VPWR VGND _08280_ sg13g2_nor3_1
X_15388_ _08040_ _08044_ _07742_ VPWR VGND _08281_ sg13g2_a21o_1
X_15389_ _07959_ _07789_ VPWR VGND _08282_ sg13g2_or2_1
X_15390_ _08037_ _08051_ _08264_ _08282_ _07741_ VPWR 
+ VGND
+ _08283_ sg13g2_a221oi_1
X_15391_ spike_o _08049_ _08253_ _08061_ VPWR VGND 
+ _08284_
+ sg13g2_and4_1
X_15392_ _07959_ _07715_ VPWR VGND _08285_ sg13g2_nand2b_1
X_15393_ spike_o _08049_ _08285_ VPWR VGND _08286_ sg13g2_a21oi_1
X_15394_ _07959_ _07936_ _07834_ _08253_ VPWR VGND 
+ _08287_
+ sg13g2_nor4_1
X_15395_ _08284_ _08286_ _08287_ VPWR VGND _08288_ sg13g2_nor3_1
X_15396_ _08256_ _08258_ _08283_ _08288_ VPWR VGND 
+ _08289_
+ sg13g2_a22oi_1
X_15397_ _08271_ _08280_ _08281_ _08289_ VPWR VGND 
+ _08290_
+ sg13g2_a22oi_1
X_15398_ _08290_ VPWR VGND _08291_ sg13g2_buf_1
X_15399_ _08022_ _08107_ VPWR VGND _08292_ sg13g2_nor2_1
X_15400_ _07755_ _08049_ _08292_ VPWR VGND _08293_ sg13g2_nand3_1
X_15401_ _08097_ _08098_ _08293_ VPWR VGND _08294_ sg13g2_and3_1
X_15402_ _07753_ _07834_ _08022_ _08292_ VPWR VGND 
+ _08295_
+ sg13g2_nor4_1
X_15403_ _08096_ _08294_ _08295_ VPWR VGND _08296_ sg13g2_a21oi_1
X_15404_ _08264_ _08094_ _08296_ VPWR VGND _08297_ sg13g2_nand3_1
X_15405_ _08264_ _08094_ _08296_ VPWR VGND _08298_ sg13g2_a21o_1
X_15406_ _08297_ _08298_ VPWR VGND _08299_ sg13g2_nand2_1
X_15407_ _07744_ _08299_ VPWR VGND _08300_ sg13g2_xnor2_1
X_15408_ _08291_ _08300_ VPWR VGND _08301_ sg13g2_xnor2_1
X_15409_ _08276_ _08301_ VPWR VGND _08302_ sg13g2_nor2_1
X_15410_ _00160_ _08276_ _08302_ VPWR VGND _08303_ sg13g2_a21oi_1
X_15411_ _07995_ _08303_ VPWR VGND _00217_ sg13g2_nor2_1
X_15412_ _08271_ _08280_ _08281_ _08289_ _07744_ VPWR 
+ VGND
+ _08304_ sg13g2_a221oi_1
X_15413_ _07744_ VPWR VGND _08305_ sg13g2_inv_1
X_15414_ _08305_ _08264_ _08094_ _08296_ VPWR VGND 
+ _08306_
+ sg13g2_and4_1
X_15415_ _07936_ _07834_ _08022_ VPWR VGND _08307_ sg13g2_nor3_1
X_15416_ _08307_ VPWR VGND _08308_ sg13g2_buf_2
X_15417_ _08107_ _08308_ VPWR VGND _08309_ sg13g2_nand2_1
X_15418_ _08096_ _08294_ VPWR VGND _08310_ sg13g2_nand2_1
X_15419_ _08264_ _08094_ _08309_ _08310_ _07744_ VPWR 
+ VGND
+ _08311_ sg13g2_a221oi_1
X_15420_ _08304_ _08306_ _08311_ VPWR VGND _08312_ sg13g2_or3_1
X_15421_ _08312_ VPWR VGND _08313_ sg13g2_buf_1
X_15422_ _08291_ _08299_ _08313_ VPWR VGND _08314_ sg13g2_a21o_1
X_15423_ _08264_ _08094_ VPWR VGND _08315_ sg13g2_nand2_1
X_15424_ _08096_ _08100_ VPWR VGND _08316_ sg13g2_nand2_1
X_15425_ spike_o _08049_ _08253_ VPWR VGND _08317_ sg13g2_nand3_1
X_15426_ _08317_ VPWR VGND _08318_ sg13g2_buf_2
X_15427_ _08318_ VPWR VGND _08319_ sg13g2_buf_8
X_15428_ _08144_ _08319_ VPWR VGND _08320_ sg13g2_nor2_1
X_15429_ _08264_ _08316_ _08139_ _08319_ _08320_ VPWR 
+ VGND
+ _08321_ sg13g2_a221oi_1
X_15430_ _08321_ VPWR VGND _08322_ sg13g2_buf_1
X_15431_ _07936_ _07834_ _08022_ _08144_ VPWR VGND 
+ _08323_
+ sg13g2_or4_1
X_15432_ _08134_ _08135_ _08319_ VPWR VGND _08324_ sg13g2_and3_1
X_15433_ _08133_ _08324_ VPWR VGND _08325_ sg13g2_nand2_1
X_15434_ _08116_ _08113_ _08323_ _08325_ _08278_ VPWR 
+ VGND
+ _08326_ sg13g2_a221oi_1
X_15435_ _08315_ _08322_ _08326_ VPWR VGND _08327_ sg13g2_a21oi_1
X_15436_ _07743_ _08327_ VPWR VGND _08328_ sg13g2_xnor2_1
X_15437_ _08314_ _08328_ VPWR VGND _08329_ sg13g2_xnor2_1
X_15438_ _00161_ _08262_ VPWR VGND _08330_ sg13g2_nor2_1
X_15439_ _08009_ _07917_ _08329_ _08262_ _08330_ VPWR 
+ VGND
+ _00218_ sg13g2_a221oi_1
X_15440_ _00162_ _08276_ VPWR VGND _08331_ sg13g2_nand2_1
X_15441_ _08297_ _08298_ _08322_ _08315_ _08326_ VPWR 
+ VGND
+ _08332_ sg13g2_a221oi_1
X_15442_ _08313_ _08327_ _08332_ _08291_ VPWR VGND 
+ _08333_
+ sg13g2_a22oi_1
X_15443_ _07775_ _08291_ VPWR VGND _08334_ sg13g2_and2_1
X_15444_ _08133_ _08324_ _08320_ VPWR VGND _08335_ sg13g2_a21oi_1
X_15445_ _08278_ _08335_ VPWR VGND _08336_ sg13g2_nor2_1
X_15446_ _08116_ _08113_ VPWR VGND _08337_ sg13g2_nand2_1
X_15447_ _08315_ _08322_ _08336_ _08337_ _07743_ VPWR 
+ VGND
+ _08338_ sg13g2_a221oi_1
X_15448_ _07775_ _08313_ _08334_ _08299_ _08338_ VPWR 
+ VGND
+ _08339_ sg13g2_a221oi_1
X_15449_ _08339_ VPWR VGND _08340_ sg13g2_buf_1
X_15450_ _08333_ _08340_ VPWR VGND _08341_ sg13g2_and2_1
X_15451_ _08162_ _08308_ VPWR VGND _08342_ sg13g2_nand2_1
X_15452_ _08165_ _08168_ _08319_ VPWR VGND _08343_ sg13g2_o21ai_1
X_15453_ _08342_ _08343_ VPWR VGND _08344_ sg13g2_nand2_1
X_15454_ _08096_ _08100_ _08133_ _08137_ VPWR VGND 
+ _08345_
+ sg13g2_nand4_1
X_15455_ _07809_ _07936_ _08345_ VPWR VGND _08346_ sg13g2_nand3_1
X_15456_ _08315_ _08344_ _08346_ VPWR VGND _08347_ sg13g2_nand3_1
X_15457_ _08347_ VPWR VGND _08348_ sg13g2_buf_1
X_15458_ _08315_ _08346_ _08344_ VPWR VGND _08349_ sg13g2_a21o_1
X_15459_ _08349_ VPWR VGND _08350_ sg13g2_buf_1
X_15460_ _08348_ _08350_ _07781_ VPWR VGND _08351_ sg13g2_a21oi_1
X_15461_ _07781_ _08348_ _08350_ VPWR VGND _08352_ sg13g2_nand3_1
X_15462_ _08352_ VPWR VGND _08353_ sg13g2_buf_1
X_15463_ _08351_ _08353_ VPWR VGND _08354_ sg13g2_nor2b_1
X_15464_ _08341_ _08354_ VPWR VGND _08355_ sg13g2_xnor2_1
X_15465_ _08262_ _08355_ VPWR VGND _08356_ sg13g2_nand2_1
X_15466_ _08331_ _08356_ _07995_ VPWR VGND _00219_ sg13g2_a21oi_1
X_15467_ _00163_ _08276_ VPWR VGND _08357_ sg13g2_nand2_1
X_15468_ _08341_ _08351_ _08353_ VPWR VGND _08358_ sg13g2_o21ai_1
X_15469_ _08195_ _08319_ VPWR VGND _08359_ sg13g2_nor2_1
X_15470_ _08198_ _08199_ _08319_ VPWR VGND _08360_ sg13g2_and3_1
X_15471_ _08360_ VPWR VGND _08361_ sg13g2_buf_4
X_15472_ _08359_ _08361_ VPWR VGND _08362_ sg13g2_or2_1
X_15473_ _08107_ _08320_ VPWR VGND _08363_ sg13g2_nand2_1
X_15474_ _08308_ _08345_ _08363_ VPWR VGND _08364_ sg13g2_o21ai_1
X_15475_ _08116_ _08342_ _08343_ VPWR VGND _08365_ sg13g2_and3_1
X_15476_ _08364_ _08365_ _08278_ VPWR VGND _08366_ sg13g2_a21oi_1
X_15477_ _08362_ _08366_ VPWR VGND _08367_ sg13g2_xnor2_1
X_15478_ _07736_ _08367_ VPWR VGND _08368_ sg13g2_xor2_1
X_15479_ _08358_ _08368_ VPWR VGND _08369_ sg13g2_xnor2_1
X_15480_ _08369_ _08262_ VPWR VGND _08370_ sg13g2_nand2b_1
X_15481_ _08357_ _08370_ _07919_ VPWR VGND _00220_ sg13g2_a21oi_1
X_15482_ _08348_ _08350_ VPWR VGND _08371_ sg13g2_nand2_1
X_15483_ _08333_ _08340_ _08371_ _07737_ _08367_ VPWR 
+ VGND
+ _08372_ sg13g2_a221oi_1
X_15484_ _07736_ _08353_ _08367_ VPWR VGND _08373_ sg13g2_a21oi_1
X_15485_ _08333_ _08340_ _08371_ _07737_ _07736_ VPWR 
+ VGND
+ _08374_ sg13g2_a221oi_1
X_15486_ _07736_ _08353_ VPWR VGND _08375_ sg13g2_nor2_1
X_15487_ _08372_ _08373_ _08374_ _08375_ VPWR VGND 
+ _08376_
+ sg13g2_or4_1
X_15488_ _08376_ VPWR VGND _08377_ sg13g2_buf_1
X_15489_ _08229_ _08319_ VPWR VGND _08378_ sg13g2_nor2_1
X_15490_ _08224_ _08319_ _08378_ VPWR VGND _08379_ sg13g2_a21o_1
X_15491_ _08379_ VPWR VGND _08380_ sg13g2_buf_1
X_15492_ _08342_ _08343_ VPWR VGND _08381_ sg13g2_and2_1
X_15493_ _08109_ _08308_ VPWR VGND _08382_ sg13g2_nand2_1
X_15494_ _08094_ _08308_ _08382_ VPWR VGND _08383_ sg13g2_o21ai_1
X_15495_ _08381_ _08364_ _08383_ _08362_ VPWR VGND 
+ _08384_
+ sg13g2_and4_1
X_15496_ _08384_ _08264_ VPWR VGND _08385_ sg13g2_nand2b_1
X_15497_ _08380_ _08385_ VPWR VGND _08386_ sg13g2_xor2_1
X_15498_ _08377_ _08386_ VPWR VGND _08387_ sg13g2_xor2_1
X_15499_ _08276_ _08387_ _07738_ VPWR VGND _08388_ sg13g2_o21ai_1
X_15500_ _07738_ _08276_ _08387_ VPWR VGND _08389_ sg13g2_or3_1
X_15501_ _08388_ _08389_ _07919_ VPWR VGND _00221_ sg13g2_a21oi_1
X_15502_ _07738_ _00092_ _08278_ VPWR VGND _08390_ sg13g2_nand3_1
X_15503_ _00092_ _08278_ _08390_ VPWR VGND _08391_ sg13g2_o21ai_1
X_15504_ _08380_ _08385_ VPWR VGND _08392_ sg13g2_nand2_1
X_15505_ _07738_ _08392_ _08262_ VPWR VGND _08393_ sg13g2_o21ai_1
X_15506_ _08386_ _08391_ _08393_ VPWR VGND _08394_ sg13g2_a21o_1
X_15507_ _08278_ _08380_ _08384_ VPWR VGND _08395_ sg13g2_nor3_1
X_15508_ _07738_ _08395_ VPWR VGND _08396_ sg13g2_xor2_1
X_15509_ _08278_ _08396_ VPWR VGND _08397_ sg13g2_nor2_1
X_15510_ _08220_ _08264_ _08392_ VPWR VGND _08398_ sg13g2_o21ai_1
X_15511_ _08397_ _08398_ _08377_ VPWR VGND _08399_ sg13g2_mux2_1
X_15512_ _07739_ _07992_ VPWR VGND _08400_ sg13g2_and2_1
X_15513_ _08394_ _08399_ _08400_ VPWR VGND _08401_ sg13g2_o21ai_1
X_15514_ _07739_ _07919_ _08394_ _08399_ VPWR VGND 
+ _08402_
+ sg13g2_or4_1
X_15515_ _08401_ _08402_ VPWR VGND _00222_ sg13g2_nand2_1
X_15516_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2635_o[0]\ VPWR VGND _08403_ sg13g2_buf_1
X_15517_ _08403_ _07799_ VPWR VGND _08404_ sg13g2_nand2_1
X_15518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[11]\ VPWR VGND _08405_ sg13g2_buf_1
X_15519_ _08405_ VPWR VGND _08406_ sg13g2_buf_2
X_15520_ _08406_ VPWR VGND _08407_ sg13g2_buf_2
X_15521_ _08407_ VPWR VGND _08408_ sg13g2_buf_2
X_15522_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[11]\ VPWR VGND _08409_ sg13g2_buf_1
X_15523_ _08409_ VPWR VGND _08410_ sg13g2_inv_1
X_15524_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[9]\ VPWR VGND _08411_ sg13g2_buf_1
X_15525_ _08411_ VPWR VGND _08412_ sg13g2_buf_1
X_15526_ _08412_ VPWR VGND _08413_ sg13g2_buf_2
X_15527_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[9]\ VPWR VGND _08414_ sg13g2_buf_1
X_15528_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[8]\ VPWR VGND _08415_ sg13g2_buf_2
X_15529_ _08415_ VPWR VGND _08416_ sg13g2_buf_4
X_15530_ _08416_ VPWR VGND _08417_ sg13g2_buf_4
X_15531_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[8]\ VPWR VGND _08418_ sg13g2_buf_1
X_15532_ _08417_ _08418_ VPWR VGND _08419_ sg13g2_nor2_1
X_15533_ _08419_ VPWR VGND _08420_ sg13g2_inv_1
X_15534_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[7]\ VPWR VGND _08421_ sg13g2_buf_2
X_15535_ _08421_ VPWR VGND _08422_ sg13g2_buf_2
X_15536_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[6]\ VPWR VGND _08423_ sg13g2_buf_2
X_15537_ _08423_ VPWR VGND _08424_ sg13g2_buf_8
X_15538_ _08424_ VPWR VGND _08425_ sg13g2_buf_4
X_15539_ _08425_ VPWR VGND _08426_ sg13g2_buf_8
X_15540_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[6]\ VPWR VGND _08427_ sg13g2_buf_1
X_15541_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[7]\ VPWR VGND _08428_ sg13g2_buf_1
X_15542_ _08426_ _08427_ _08428_ VPWR VGND _08429_ sg13g2_a21o_1
X_15543_ _08426_ _08428_ _08427_ VPWR VGND _08430_ sg13g2_and3_1
X_15544_ _08422_ _08429_ _08430_ VPWR VGND _08431_ sg13g2_a21o_1
X_15545_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[10]\ VPWR VGND _08432_ sg13g2_buf_2
X_15546_ _08432_ VPWR VGND _08433_ sg13g2_buf_2
X_15547_ _08433_ VPWR VGND _08434_ sg13g2_buf_2
X_15548_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[10]\ VPWR VGND _08435_ sg13g2_buf_1
X_15549_ _08416_ VPWR VGND _08436_ sg13g2_buf_2
X_15550_ _08434_ _08435_ _08418_ _08436_ VPWR VGND 
+ _08437_
+ sg13g2_a22oi_1
X_15551_ _08437_ VPWR VGND _08438_ sg13g2_inv_1
X_15552_ _08413_ _08414_ _08420_ _08431_ _08438_ VPWR 
+ VGND
+ _08439_ sg13g2_a221oi_1
X_15553_ _08439_ VPWR VGND _08440_ sg13g2_buf_2
X_15554_ _08433_ VPWR VGND _08441_ sg13g2_buf_2
X_15555_ _08411_ VPWR VGND _08442_ sg13g2_inv_1
X_15556_ _08442_ VPWR VGND _08443_ sg13g2_buf_1
X_15557_ _08414_ VPWR VGND _08444_ sg13g2_inv_1
X_15558_ _08434_ _08435_ VPWR VGND _08445_ sg13g2_nand2_1
X_15559_ _08443_ _08444_ _08445_ VPWR VGND _08446_ sg13g2_nand3_1
X_15560_ _08441_ _08435_ _08446_ VPWR VGND _08447_ sg13g2_o21ai_1
X_15561_ _08447_ VPWR VGND _08448_ sg13g2_buf_1
X_15562_ _08410_ _08440_ _08448_ VPWR VGND _08449_ sg13g2_nor3_1
X_15563_ _08440_ _08448_ _08410_ VPWR VGND _08450_ sg13g2_o21ai_1
X_15564_ _08408_ _08449_ _08450_ VPWR VGND _08451_ sg13g2_o21ai_1
X_15565_ _08451_ VPWR VGND _08452_ sg13g2_buf_2
X_15566_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[12]\ VPWR VGND _08453_ sg13g2_buf_1
X_15567_ _08453_ VPWR VGND _08454_ sg13g2_buf_2
X_15568_ _08454_ VPWR VGND _08455_ sg13g2_buf_1
X_15569_ _08455_ VPWR VGND _08456_ sg13g2_buf_2
X_15570_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[12]\ VPWR VGND _08457_ sg13g2_buf_1
X_15571_ _08456_ _08457_ VPWR VGND _08458_ sg13g2_nand2_1
X_15572_ _08456_ _08457_ VPWR VGND _08459_ sg13g2_nor2_1
X_15573_ _08452_ _08458_ _08459_ VPWR VGND _08460_ sg13g2_a21oi_1
X_15574_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[13]\ VPWR VGND _08461_ sg13g2_buf_1
X_15575_ _08461_ VPWR VGND _08462_ sg13g2_buf_1
X_15576_ _08462_ VPWR VGND _08463_ sg13g2_buf_1
X_15577_ _08463_ VPWR VGND _08464_ sg13g2_buf_1
X_15578_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[13]\ VPWR VGND _08465_ sg13g2_buf_1
X_15579_ _08464_ _08465_ VPWR VGND _08466_ sg13g2_xor2_1
X_15580_ _08460_ _08466_ VPWR VGND _08467_ sg13g2_xnor2_1
X_15581_ _00067_ VPWR VGND _08468_ sg13g2_buf_1
X_15582_ _08422_ VPWR VGND _08469_ sg13g2_buf_2
X_15583_ _08469_ _08428_ VPWR VGND _08470_ sg13g2_xor2_1
X_15584_ _08468_ _08470_ VPWR VGND _08471_ sg13g2_and2_1
X_15585_ _08471_ VPWR VGND _08472_ sg13g2_buf_1
X_15586_ _00068_ VPWR VGND _08473_ sg13g2_buf_1
X_15587_ _08473_ VPWR VGND _08474_ sg13g2_buf_1
X_15588_ _08474_ VPWR VGND _08475_ sg13g2_inv_1
X_15589_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[5]\ VPWR VGND _08476_ sg13g2_buf_1
X_15590_ _08476_ VPWR VGND _08477_ sg13g2_inv_1
X_15591_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ VPWR VGND _08478_ sg13g2_buf_1
X_15592_ _08477_ _08478_ VPWR VGND _08479_ sg13g2_nor2_1
X_15593_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[4]\ VPWR VGND _08480_ sg13g2_buf_1
X_15594_ _08480_ VPWR VGND _08481_ sg13g2_inv_1
X_15595_ _08481_ VPWR VGND _08482_ sg13g2_buf_1
X_15596_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[4]\ VPWR VGND _08483_ sg13g2_buf_1
X_15597_ _08482_ _08483_ VPWR VGND _08484_ sg13g2_nand2_1
X_15598_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[3]\ VPWR VGND _08485_ sg13g2_buf_1
X_15599_ _08485_ VPWR VGND _08486_ sg13g2_inv_1
X_15600_ _08486_ VPWR VGND _08487_ sg13g2_buf_1
X_15601_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ VPWR VGND _08488_ sg13g2_inv_1
X_15602_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[2]\ VPWR VGND _08489_ sg13g2_buf_1
X_15603_ _08489_ VPWR VGND _08490_ sg13g2_inv_1
X_15604_ _08490_ VPWR VGND _08491_ sg13g2_buf_1
X_15605_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[2]\ VPWR VGND _08492_ sg13g2_buf_1
X_15606_ _08491_ _08492_ VPWR VGND _08493_ sg13g2_nor2_1
X_15607_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[0]\ VPWR VGND _08494_ sg13g2_buf_1
X_15608_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ VPWR VGND _08495_ sg13g2_buf_1
X_15609_ _08494_ _08495_ VPWR VGND _08496_ sg13g2_nor2b_1
X_15610_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ VPWR VGND _08497_ sg13g2_buf_1
X_15611_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[1]\ VPWR VGND _08498_ sg13g2_buf_2
X_15612_ _08497_ _08498_ VPWR VGND _08499_ sg13g2_nand2b_1
X_15613_ _08498_ _08497_ VPWR VGND _08500_ sg13g2_nor2b_1
X_15614_ _08491_ _08492_ _08496_ _08499_ _08500_ VPWR 
+ VGND
+ _08501_ sg13g2_a221oi_1
X_15615_ _08488_ _08493_ _08501_ VPWR VGND _08502_ sg13g2_nor3_1
X_15616_ _08493_ _08501_ _08488_ VPWR VGND _08503_ sg13g2_o21ai_1
X_15617_ _08487_ _08502_ _08503_ VPWR VGND _08504_ sg13g2_o21ai_1
X_15618_ _08482_ _08483_ VPWR VGND _08505_ sg13g2_nor2_1
X_15619_ _08484_ _08504_ _08505_ VPWR VGND _08506_ sg13g2_a21o_1
X_15620_ _08506_ VPWR VGND _08507_ sg13g2_buf_1
X_15621_ _08474_ VPWR VGND _08508_ sg13g2_buf_1
X_15622_ _08476_ _08478_ VPWR VGND _08509_ sg13g2_nor2b_1
X_15623_ _08508_ _08509_ VPWR VGND _08510_ sg13g2_nor2_1
X_15624_ _08427_ VPWR VGND _08511_ sg13g2_inv_1
X_15625_ _08475_ _08479_ _08507_ _08510_ _08511_ VPWR 
+ VGND
+ _08512_ sg13g2_a221oi_1
X_15626_ _08426_ VPWR VGND _08513_ sg13g2_buf_1
X_15627_ _08513_ VPWR VGND _08514_ sg13g2_buf_2
X_15628_ _08514_ VPWR VGND _08515_ sg13g2_inv_1
X_15629_ _08515_ VPWR VGND _08516_ sg13g2_buf_1
X_15630_ _08485_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ VPWR VGND _08517_ sg13g2_xor2_1
X_15631_ _08494_ VPWR VGND _08518_ sg13g2_buf_2
X_15632_ _08518_ _08495_ VPWR VGND _08519_ sg13g2_xnor2_1
X_15633_ _08480_ _08483_ VPWR VGND _08520_ sg13g2_xnor2_1
X_15634_ _08489_ _08492_ VPWR VGND _08521_ sg13g2_xnor2_1
X_15635_ _08498_ _08497_ VPWR VGND _08522_ sg13g2_xnor2_1
X_15636_ _08519_ _08520_ _08521_ _08522_ VPWR VGND 
+ _08523_
+ sg13g2_nand4_1
X_15637_ _08479_ _08509_ _08517_ _08523_ VPWR VGND 
+ _08524_
+ sg13g2_nor4_1
X_15638_ _08474_ _08427_ VPWR VGND _08525_ sg13g2_xnor2_1
X_15639_ _08525_ _08472_ VPWR VGND _08526_ sg13g2_nor2_1
X_15640_ _08468_ VPWR VGND _08527_ sg13g2_buf_1
X_15641_ _08527_ _08470_ VPWR VGND _08528_ sg13g2_nor2_1
X_15642_ _08524_ _08526_ _08528_ VPWR VGND _08529_ sg13g2_a21oi_1
X_15643_ _08516_ _08529_ VPWR VGND _08530_ sg13g2_and2_1
X_15644_ _08472_ _08512_ _08530_ VPWR VGND _08531_ sg13g2_o21ai_1
X_15645_ _08468_ VPWR VGND _08532_ sg13g2_inv_1
X_15646_ _08532_ VPWR VGND _08533_ sg13g2_buf_1
X_15647_ _08533_ VPWR VGND _08534_ sg13g2_buf_1
X_15648_ _08534_ _08511_ _08470_ VPWR VGND _08535_ sg13g2_nor3_1
X_15649_ _08475_ _08479_ _08507_ _08510_ _08427_ VPWR 
+ VGND
+ _08536_ sg13g2_a221oi_1
X_15650_ _08427_ _08470_ VPWR VGND _08537_ sg13g2_and2_1
X_15651_ _08474_ _08427_ _08470_ VPWR VGND _08538_ sg13g2_nor3_1
X_15652_ _08533_ _08525_ _08537_ _08508_ _08538_ VPWR 
+ VGND
+ _08539_ sg13g2_a221oi_1
X_15653_ _08539_ _08524_ VPWR VGND _08540_ sg13g2_nor2b_1
X_15654_ _08534_ _08537_ _08540_ VPWR VGND _08541_ sg13g2_a21o_1
X_15655_ _08514_ VPWR VGND _08542_ sg13g2_buf_2
X_15656_ _08542_ VPWR VGND _08543_ sg13g2_buf_2
X_15657_ _08511_ _08528_ VPWR VGND _08544_ sg13g2_nand2_1
X_15658_ _08543_ _08529_ _08544_ VPWR VGND _08545_ sg13g2_o21ai_1
X_15659_ _08516_ _08541_ _08545_ VPWR VGND _08546_ sg13g2_nor3_1
X_15660_ _08535_ _08536_ _08546_ VPWR VGND _08547_ sg13g2_o21ai_1
X_15661_ _00076_ VPWR VGND _08548_ sg13g2_buf_1
X_15662_ _08548_ VPWR VGND _08549_ sg13g2_buf_1
X_15663_ _08436_ VPWR VGND _08550_ sg13g2_buf_2
X_15664_ _08550_ VPWR VGND _08551_ sg13g2_buf_2
X_15665_ _08551_ _08418_ VPWR VGND _08552_ sg13g2_xor2_1
X_15666_ _08431_ _08552_ VPWR VGND _08553_ sg13g2_xnor2_1
X_15667_ _08549_ _08553_ VPWR VGND _08554_ sg13g2_xnor2_1
X_15668_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[6]\ VPWR VGND _08555_ sg13g2_buf_1
X_15669_ _08555_ VPWR VGND _08556_ sg13g2_buf_1
X_15670_ _08556_ VPWR VGND _08557_ sg13g2_buf_1
X_15671_ _08557_ _08479_ _08507_ VPWR VGND _08558_ sg13g2_nor3_1
X_15672_ _08513_ _08473_ VPWR VGND _08559_ sg13g2_xor2_1
X_15673_ _08559_ VPWR VGND _08560_ sg13g2_buf_1
X_15674_ _08427_ _08560_ _08509_ VPWR VGND _08561_ sg13g2_a21oi_1
X_15675_ _08557_ _08560_ VPWR VGND _08562_ sg13g2_nor2_1
X_15676_ _08472_ _08562_ _08511_ VPWR VGND _08563_ sg13g2_o21ai_1
X_15677_ _08557_ _08561_ _08563_ VPWR VGND _08564_ sg13g2_o21ai_1
X_15678_ _08543_ _08541_ _08545_ VPWR VGND _08565_ sg13g2_a21oi_1
X_15679_ _08558_ _08564_ _08565_ VPWR VGND _08566_ sg13g2_o21ai_1
X_15680_ _08531_ _08547_ _08554_ _08566_ VPWR VGND 
+ _08567_
+ sg13g2_nand4_1
X_15681_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[12]\ VPWR VGND _08568_ sg13g2_buf_1
X_15682_ _08568_ VPWR VGND _08569_ sg13g2_inv_1
X_15683_ _08456_ VPWR VGND _08570_ sg13g2_buf_1
X_15684_ _08570_ _08457_ VPWR VGND _08571_ sg13g2_xor2_1
X_15685_ _08452_ _08571_ VPWR VGND _08572_ sg13g2_xnor2_1
X_15686_ _08569_ _08572_ VPWR VGND _08573_ sg13g2_nor2_1
X_15687_ _00075_ VPWR VGND _08574_ sg13g2_buf_1
X_15688_ _08574_ VPWR VGND _08575_ sg13g2_buf_1
X_15689_ _08575_ VPWR VGND _08576_ sg13g2_buf_1
X_15690_ _08576_ VPWR VGND _08577_ sg13g2_buf_1
X_15691_ _08469_ VPWR VGND _08578_ sg13g2_buf_2
X_15692_ _08436_ _08418_ _08429_ _08578_ _08430_ VPWR 
+ VGND
+ _08579_ sg13g2_a221oi_1
X_15693_ _08579_ VPWR VGND _08580_ sg13g2_buf_1
X_15694_ _08419_ _08580_ VPWR VGND _08581_ sg13g2_nor2_1
X_15695_ _08413_ VPWR VGND _08582_ sg13g2_buf_2
X_15696_ _08582_ VPWR VGND _08583_ sg13g2_buf_2
X_15697_ _08583_ VPWR VGND _08584_ sg13g2_buf_2
X_15698_ _08584_ _08414_ VPWR VGND _08585_ sg13g2_xnor2_1
X_15699_ _08581_ _08585_ VPWR VGND _08586_ sg13g2_xnor2_1
X_15700_ _08577_ _08586_ VPWR VGND _08587_ sg13g2_nor2_1
X_15701_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[10]\ VPWR VGND _08588_ sg13g2_buf_1
X_15702_ _08588_ VPWR VGND _08589_ sg13g2_buf_1
X_15703_ _08583_ VPWR VGND _08590_ sg13g2_buf_1
X_15704_ _08444_ _08419_ _08580_ VPWR VGND _08591_ sg13g2_nor3_1
X_15705_ _08419_ _08580_ _08444_ VPWR VGND _08592_ sg13g2_o21ai_1
X_15706_ _08590_ _08591_ _08592_ VPWR VGND _08593_ sg13g2_o21ai_1
X_15707_ _08441_ VPWR VGND _08594_ sg13g2_buf_2
X_15708_ _08594_ VPWR VGND _08595_ sg13g2_buf_1
X_15709_ _08595_ _08435_ VPWR VGND _08596_ sg13g2_xnor2_1
X_15710_ _08593_ _08596_ VPWR VGND _08597_ sg13g2_xnor2_1
X_15711_ _08440_ _08448_ VPWR VGND _08598_ sg13g2_nor2_1
X_15712_ _08408_ _08409_ VPWR VGND _08599_ sg13g2_xnor2_1
X_15713_ _08598_ _08599_ VPWR VGND _08600_ sg13g2_xor2_1
X_15714_ _00073_ VPWR VGND _08601_ sg13g2_buf_1
X_15715_ _08601_ VPWR VGND _08602_ sg13g2_inv_1
X_15716_ _08589_ _08597_ _08600_ _08602_ VPWR VGND 
+ _08603_
+ sg13g2_a22oi_1
X_15717_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[8]\ VPWR VGND _08604_ sg13g2_buf_1
X_15718_ _08604_ VPWR VGND _08605_ sg13g2_buf_1
X_15719_ _08605_ _08553_ VPWR VGND _08606_ sg13g2_nand2_1
X_15720_ _08587_ _08603_ _08606_ VPWR VGND _08607_ sg13g2_nand3b_1
X_15721_ _08573_ _08607_ VPWR VGND _08608_ sg13g2_nor2_1
X_15722_ _08454_ VPWR VGND _08609_ sg13g2_buf_1
X_15723_ _00072_ VPWR VGND _08610_ sg13g2_buf_1
X_15724_ _08609_ _08610_ VPWR VGND _08611_ sg13g2_xnor2_1
X_15725_ _08611_ VPWR VGND _08612_ sg13g2_buf_1
X_15726_ _08457_ _08612_ VPWR VGND _08613_ sg13g2_xor2_1
X_15727_ _08440_ _08448_ _08599_ VPWR VGND _08614_ sg13g2_nor3_1
X_15728_ _08601_ VPWR VGND _08615_ sg13g2_buf_1
X_15729_ _08408_ VPWR VGND _08616_ sg13g2_buf_1
X_15730_ _08616_ VPWR VGND _08617_ sg13g2_buf_1
X_15731_ _08617_ _08409_ VPWR VGND _08618_ sg13g2_nand2_1
X_15732_ _08615_ _08598_ _08618_ VPWR VGND _08619_ sg13g2_a21oi_1
X_15733_ _08614_ _08619_ VPWR VGND _08620_ sg13g2_nor2_1
X_15734_ _08441_ _00074_ VPWR VGND _08621_ sg13g2_xnor2_1
X_15735_ _08621_ VPWR VGND _08622_ sg13g2_buf_1
X_15736_ _08622_ VPWR VGND _08623_ sg13g2_buf_1
X_15737_ _08435_ _08623_ VPWR VGND _08624_ sg13g2_xnor2_1
X_15738_ _08443_ VPWR VGND _08625_ sg13g2_buf_1
X_15739_ _08576_ VPWR VGND _08626_ sg13g2_buf_1
X_15740_ _08626_ _08591_ _08592_ VPWR VGND _08627_ sg13g2_o21ai_1
X_15741_ _08626_ _08592_ VPWR VGND _08628_ sg13g2_nor2_1
X_15742_ _08625_ _08627_ _08628_ VPWR VGND _08629_ sg13g2_a21oi_1
X_15743_ _08419_ _08580_ _08585_ VPWR VGND _08630_ sg13g2_nor3_1
X_15744_ _08590_ _08414_ VPWR VGND _08631_ sg13g2_nand2_1
X_15745_ _08626_ _08581_ _08631_ VPWR VGND _08632_ sg13g2_a21oi_1
X_15746_ _08630_ _08632_ _08624_ VPWR VGND _08633_ sg13g2_nor3_1
X_15747_ _08624_ _08629_ _08633_ VPWR VGND _08634_ sg13g2_a21o_1
X_15748_ _08602_ VPWR VGND _08635_ sg13g2_buf_1
X_15749_ _08409_ _08598_ VPWR VGND _08636_ sg13g2_nor2_1
X_15750_ _08601_ _08449_ _08450_ VPWR VGND _08637_ sg13g2_o21ai_1
X_15751_ _08406_ VPWR VGND _08638_ sg13g2_inv_1
X_15752_ _08638_ VPWR VGND _08639_ sg13g2_buf_1
X_15753_ _08635_ _08636_ _08637_ _08639_ _08613_ VPWR 
+ VGND
+ _08640_ sg13g2_a221oi_1
X_15754_ _08613_ _08620_ _08634_ _08603_ _08640_ VPWR 
+ VGND
+ _08641_ sg13g2_a221oi_1
X_15755_ _08573_ _08641_ VPWR VGND _08642_ sg13g2_nor2_1
X_15756_ _08567_ _08608_ _08642_ VPWR VGND _08643_ sg13g2_a21oi_1
X_15757_ _00071_ VPWR VGND _08644_ sg13g2_buf_1
X_15758_ _08644_ VPWR VGND _08645_ sg13g2_inv_1
X_15759_ _08645_ VPWR VGND _08646_ sg13g2_buf_1
X_15760_ _08467_ _08643_ _08646_ VPWR VGND _08647_ sg13g2_o21ai_1
X_15761_ _08467_ _08643_ VPWR VGND _08648_ sg13g2_nand2_1
X_15762_ _08647_ _08648_ VPWR VGND _08649_ sg13g2_nand2_1
X_15763_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[14]\ VPWR VGND _08650_ sg13g2_buf_1
X_15764_ _08650_ VPWR VGND _08651_ sg13g2_buf_1
X_15765_ _08651_ VPWR VGND _08652_ sg13g2_buf_1
X_15766_ _08652_ VPWR VGND _08653_ sg13g2_buf_1
X_15767_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[14]\ VPWR VGND _08654_ sg13g2_buf_1
X_15768_ _08653_ _08654_ VPWR VGND _08655_ sg13g2_and2_1
X_15769_ _08654_ _08465_ VPWR VGND _08656_ sg13g2_nand2_1
X_15770_ _08652_ _08465_ VPWR VGND _08657_ sg13g2_nand2_1
X_15771_ _08452_ _08458_ _08656_ _08657_ _08459_ VPWR 
+ VGND
+ _08658_ sg13g2_a221oi_1
X_15772_ _08463_ _08654_ VPWR VGND _08659_ sg13g2_nand2_1
X_15773_ _08462_ VPWR VGND _08660_ sg13g2_buf_1
X_15774_ _08652_ _08660_ VPWR VGND _08661_ sg13g2_nand2_1
X_15775_ _08452_ _08458_ _08659_ _08661_ _08459_ VPWR 
+ VGND
+ _08662_ sg13g2_a221oi_1
X_15776_ _08465_ VPWR VGND _08663_ sg13g2_inv_1
X_15777_ _08659_ _08661_ _08663_ VPWR VGND _08664_ sg13g2_a21oi_1
X_15778_ _08655_ _08658_ _08662_ _08664_ VPWR VGND 
+ _08665_
+ sg13g2_nor4_1
X_15779_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[15]\ VPWR VGND _08666_ sg13g2_buf_1
X_15780_ _08666_ VPWR VGND _08667_ sg13g2_buf_1
X_15781_ _08667_ VPWR VGND _08668_ sg13g2_buf_1
X_15782_ _08668_ VPWR VGND _08669_ sg13g2_buf_1
X_15783_ _08669_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[15]\ VPWR VGND _08670_ sg13g2_xor2_1
X_15784_ _08665_ _08670_ VPWR VGND _08671_ sg13g2_xnor2_1
X_15785_ _08465_ _08460_ _08464_ VPWR VGND _08672_ sg13g2_a21o_1
X_15786_ _08465_ _08460_ _08672_ VPWR VGND _08673_ sg13g2_o21ai_1
X_15787_ _08654_ _08673_ VPWR VGND _08674_ sg13g2_xor2_1
X_15788_ _00070_ VPWR VGND _08675_ sg13g2_buf_1
X_15789_ _08650_ _08675_ VPWR VGND _08676_ sg13g2_xnor2_1
X_15790_ _08674_ _08676_ VPWR VGND _08677_ sg13g2_xnor2_1
X_15791_ _08671_ _08677_ VPWR VGND _08678_ sg13g2_nor2_1
X_15792_ _00069_ VPWR VGND _08679_ sg13g2_buf_1
X_15793_ _08679_ VPWR VGND _08680_ sg13g2_buf_1
X_15794_ _08680_ VPWR VGND _08681_ sg13g2_buf_1
X_15795_ _08653_ VPWR VGND _08682_ sg13g2_buf_1
X_15796_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[14]\ VPWR VGND _08683_ sg13g2_buf_1
X_15797_ _08683_ VPWR VGND _08684_ sg13g2_buf_1
X_15798_ _08682_ _08684_ VPWR VGND _08685_ sg13g2_nand2_1
X_15799_ _08651_ VPWR VGND _08686_ sg13g2_inv_1
X_15800_ _08686_ _08684_ VPWR VGND _08687_ sg13g2_nand2_1
X_15801_ _08685_ _08687_ _08674_ VPWR VGND _08688_ sg13g2_mux2_1
X_15802_ _08681_ _08671_ _08688_ VPWR VGND _08689_ sg13g2_a21oi_1
X_15803_ _08649_ _08678_ _08689_ VPWR VGND _08690_ sg13g2_a21oi_1
X_15804_ _08680_ _08677_ VPWR VGND _08691_ sg13g2_nor2_1
X_15805_ _08681_ _08671_ VPWR VGND _08692_ sg13g2_nor2_1
X_15806_ _08649_ _08691_ _08692_ VPWR VGND _08693_ sg13g2_a21oi_1
X_15807_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[15]\ VPWR VGND _08694_ sg13g2_inv_1
X_15808_ _08666_ VPWR VGND _08695_ sg13g2_inv_1
X_15809_ _08695_ VPWR VGND _08696_ sg13g2_buf_1
X_15810_ _08694_ _08665_ _08696_ VPWR VGND _08697_ sg13g2_o21ai_1
X_15811_ _08694_ _08665_ VPWR VGND _08698_ sg13g2_nand2_1
X_15812_ _08697_ _08698_ VPWR VGND _08699_ sg13g2_nand2_1
X_15813_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[16]\ _08699_ VPWR VGND _08700_ sg13g2_xnor2_1
X_15814_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[16]\ VPWR VGND _08701_ sg13g2_buf_1
X_15815_ _00078_ VPWR VGND _08702_ sg13g2_buf_1
X_15816_ _08701_ _08702_ VPWR VGND _08703_ sg13g2_xnor2_1
X_15817_ _08703_ VPWR VGND _08704_ sg13g2_buf_1
X_15818_ _08700_ _08704_ VPWR VGND _08705_ sg13g2_xor2_1
X_15819_ _08690_ _08693_ _08705_ VPWR VGND _08706_ sg13g2_a21oi_1
X_15820_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[17]\ VPWR VGND _08707_ sg13g2_buf_1
X_15821_ _08707_ VPWR VGND _08708_ sg13g2_buf_1
X_15822_ _08708_ VPWR VGND _08709_ sg13g2_buf_1
X_15823_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[17]\ VPWR VGND _08710_ sg13g2_buf_1
X_15824_ _08710_ VPWR VGND _08711_ sg13g2_inv_1
X_15825_ _08711_ VPWR VGND _08712_ sg13g2_buf_1
X_15826_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[17]\ VPWR VGND _08713_ sg13g2_buf_1
X_15827_ _08713_ VPWR VGND _08714_ sg13g2_inv_1
X_15828_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[16]\ VPWR VGND _08715_ sg13g2_inv_1
X_15829_ _08701_ VPWR VGND _08716_ sg13g2_inv_1
X_15830_ _08696_ _08694_ _08715_ _08716_ _08665_ VPWR 
+ VGND
+ _08717_ sg13g2_a221oi_1
X_15831_ _08716_ _08715_ VPWR VGND _08718_ sg13g2_nand2_1
X_15832_ _08668_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[15]\ _08718_ VPWR VGND _08719_ sg13g2_nand3_1
X_15833_ _08716_ _08715_ _08719_ VPWR VGND _08720_ sg13g2_o21ai_1
X_15834_ _08717_ _08720_ VPWR VGND _08721_ sg13g2_nor2_1
X_15835_ _08714_ _08721_ VPWR VGND _08722_ sg13g2_xnor2_1
X_15836_ _08712_ _08722_ VPWR VGND _08723_ sg13g2_xnor2_1
X_15837_ _08701_ VPWR VGND _08724_ sg13g2_buf_1
X_15838_ _08724_ VPWR VGND _08725_ sg13g2_buf_1
X_15839_ _08725_ VPWR VGND _08726_ sg13g2_buf_1
X_15840_ _08726_ _08700_ VPWR VGND _08727_ sg13g2_xnor2_1
X_15841_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[16]\ VPWR VGND _08728_ sg13g2_buf_1
X_15842_ _08728_ VPWR VGND _08729_ sg13g2_buf_1
X_15843_ _08709_ _08723_ _08727_ _08729_ VPWR VGND 
+ _08730_
+ sg13g2_a22oi_1
X_15844_ _08706_ _08730_ VPWR VGND _08731_ sg13g2_nand2b_1
X_15845_ _08721_ VPWR VGND _08732_ sg13g2_inv_1
X_15846_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2637_o\ VPWR VGND _08733_ sg13g2_buf_1
X_15847_ _08707_ _08733_ VPWR VGND _08734_ sg13g2_nand2_1
X_15848_ _08713_ _08734_ VPWR VGND _08735_ sg13g2_and2_1
X_15849_ _08707_ _08713_ _08732_ VPWR VGND _08736_ sg13g2_nor3_1
X_15850_ _08732_ _08735_ _08736_ VPWR VGND _08737_ sg13g2_a21oi_1
X_15851_ _08710_ VPWR VGND _08738_ sg13g2_buf_1
X_15852_ _08738_ VPWR VGND _08739_ sg13g2_buf_1
X_15853_ _08739_ VPWR VGND _08740_ sg13g2_buf_1
X_15854_ _00077_ VPWR VGND _08741_ sg13g2_buf_1
X_15855_ _08741_ VPWR VGND _08742_ sg13g2_buf_1
X_15856_ _08740_ _08734_ _08742_ VPWR VGND _08743_ sg13g2_a21oi_1
X_15857_ _08741_ VPWR VGND _08744_ sg13g2_inv_1
X_15858_ _08711_ _08744_ VPWR VGND _08745_ sg13g2_nor2_1
X_15859_ _08714_ _08733_ _08745_ VPWR VGND _08746_ sg13g2_nand3_1
X_15860_ _08713_ _08733_ _08745_ VPWR VGND _08747_ sg13g2_nand3_1
X_15861_ _08746_ _08747_ _08721_ VPWR VGND _08748_ sg13g2_mux2_1
X_15862_ _08710_ _08741_ VPWR VGND _08749_ sg13g2_xor2_1
X_15863_ _08749_ VPWR VGND _08750_ sg13g2_buf_1
X_15864_ _08713_ _08733_ _08732_ _08750_ VPWR VGND 
+ _08751_
+ sg13g2_nand4_1
X_15865_ _08714_ _08721_ _08750_ VPWR VGND _08752_ sg13g2_nand3_1
X_15866_ _08748_ _08751_ _08752_ VPWR VGND _08753_ sg13g2_nand3_1
X_15867_ _08737_ _08743_ _08753_ VPWR VGND _08754_ sg13g2_a21oi_1
X_15868_ _07733_ _08754_ VPWR VGND _08755_ sg13g2_nor2_1
X_15869_ _07795_ _08404_ _08731_ _08755_ VPWR VGND 
+ _00493_
+ sg13g2_a22oi_1
X_15870_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2647_o[0]\ VPWR VGND _08756_ sg13g2_buf_1
X_15871_ _07801_ VPWR VGND _08757_ sg13g2_inv_1
X_15872_ _08757_ VPWR VGND _08758_ sg13g2_buf_1
X_15873_ _08758_ VPWR VGND _08759_ sg13g2_buf_1
X_15874_ _08759_ VPWR VGND _08760_ sg13g2_buf_1
X_15875_ _08756_ _08760_ VPWR VGND _08761_ sg13g2_nand2_1
X_15876_ _08708_ VPWR VGND _08762_ sg13g2_inv_1
X_15877_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[16]\ VPWR VGND _08763_ sg13g2_buf_1
X_15878_ _08763_ VPWR VGND _08764_ sg13g2_inv_1
X_15879_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[13]\ VPWR VGND _08765_ sg13g2_buf_1
X_15880_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[12]\ VPWR VGND _08766_ sg13g2_buf_1
X_15881_ _08766_ VPWR VGND _08767_ sg13g2_inv_1
X_15882_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[10]\ VPWR VGND _08768_ sg13g2_buf_1
X_15883_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[8]\ VPWR VGND _08769_ sg13g2_buf_1
X_15884_ _08415_ _08769_ VPWR VGND _08770_ sg13g2_nor2_1
X_15885_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[6]\ VPWR VGND _08771_ sg13g2_buf_1
X_15886_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[7]\ VPWR VGND _08772_ sg13g2_buf_1
X_15887_ _08423_ _08771_ _08772_ VPWR VGND _08773_ sg13g2_a21o_1
X_15888_ _08423_ _08772_ _08771_ VPWR VGND _08774_ sg13g2_and3_1
X_15889_ _08415_ _08769_ _08773_ _08421_ _08774_ VPWR 
+ VGND
+ _08775_ sg13g2_a221oi_1
X_15890_ _08775_ VPWR VGND _08776_ sg13g2_buf_1
X_15891_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[9]\ VPWR VGND _08777_ sg13g2_inv_1
X_15892_ _08770_ _08776_ _08777_ VPWR VGND _08778_ sg13g2_o21ai_1
X_15893_ _08777_ _08770_ _08776_ VPWR VGND _08779_ sg13g2_nor3_1
X_15894_ _08434_ _08768_ _08778_ _08412_ _08779_ VPWR 
+ VGND
+ _08780_ sg13g2_a221oi_1
X_15895_ _08780_ VPWR VGND _08781_ sg13g2_buf_1
X_15896_ _08434_ _08768_ VPWR VGND _08782_ sg13g2_nor2_1
X_15897_ _08782_ VPWR VGND _08783_ sg13g2_buf_1
X_15898_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[11]\ VPWR VGND _08784_ sg13g2_buf_1
X_15899_ _08405_ _08784_ VPWR VGND _08785_ sg13g2_nor2_1
X_15900_ _08767_ _08781_ _08783_ _08785_ VPWR VGND 
+ _08786_
+ sg13g2_nor4_1
X_15901_ _08453_ VPWR VGND _08787_ sg13g2_inv_1
X_15902_ _08787_ _08781_ _08783_ _08785_ VPWR VGND 
+ _08788_
+ sg13g2_nor4_1
X_15903_ _08405_ _08784_ VPWR VGND _08789_ sg13g2_and2_1
X_15904_ _08453_ _08766_ _08789_ VPWR VGND _08790_ sg13g2_o21ai_1
X_15905_ _08787_ _08767_ _08790_ VPWR VGND _08791_ sg13g2_o21ai_1
X_15906_ _08765_ _08786_ _08788_ _08791_ VPWR VGND 
+ _08792_
+ sg13g2_or4_1
X_15907_ _08792_ VPWR VGND _08793_ sg13g2_buf_1
X_15908_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[15]\ VPWR VGND _08794_ sg13g2_buf_1
X_15909_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[14]\ VPWR VGND _08795_ sg13g2_buf_1
X_15910_ _08651_ _08795_ VPWR VGND _08796_ sg13g2_nand2_1
X_15911_ _08794_ _08796_ VPWR VGND _08797_ sg13g2_nand2b_1
X_15912_ _08695_ _08796_ VPWR VGND _08798_ sg13g2_nand2_1
X_15913_ _08765_ _08766_ VPWR VGND _08799_ sg13g2_nand2_1
X_15914_ _08781_ _08783_ _08785_ _08799_ VPWR VGND 
+ _08800_
+ sg13g2_nor4_1
X_15915_ _08453_ _08765_ VPWR VGND _08801_ sg13g2_nand2_1
X_15916_ _08781_ _08783_ _08785_ _08801_ VPWR VGND 
+ _08802_
+ sg13g2_nor4_1
X_15917_ _08406_ _08784_ VPWR VGND _08803_ sg13g2_nand2_1
X_15918_ _08799_ _08801_ _08803_ VPWR VGND _08804_ sg13g2_a21oi_1
X_15919_ _08767_ _08801_ VPWR VGND _08805_ sg13g2_nor2_1
X_15920_ _08800_ _08802_ _08804_ _08805_ VPWR VGND 
+ _08806_
+ sg13g2_or4_1
X_15921_ _08806_ VPWR VGND _08807_ sg13g2_buf_1
X_15922_ _08660_ _08793_ _08797_ _08798_ _08807_ VPWR 
+ VGND
+ _08808_ sg13g2_a221oi_1
X_15923_ _08808_ VPWR VGND _08809_ sg13g2_buf_1
X_15924_ _08651_ _08795_ VPWR VGND _08810_ sg13g2_or2_1
X_15925_ _08810_ VPWR VGND _08811_ sg13g2_buf_1
X_15926_ _08666_ _08794_ _08811_ VPWR VGND _08812_ sg13g2_a21o_1
X_15927_ _08666_ _08794_ _08812_ VPWR VGND _08813_ sg13g2_o21ai_1
X_15928_ _08764_ _08809_ _08813_ VPWR VGND _08814_ sg13g2_nor3_1
X_15929_ _08809_ _08813_ _08764_ VPWR VGND _08815_ sg13g2_o21ai_1
X_15930_ _08724_ _08814_ _08815_ VPWR VGND _08816_ sg13g2_o21ai_1
X_15931_ _08816_ VPWR VGND _08817_ sg13g2_buf_1
X_15932_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[17]\ _08817_ VPWR VGND _08818_ sg13g2_xnor2_1
X_15933_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[17]\ VPWR VGND _08819_ sg13g2_inv_1
X_15934_ _08738_ _08819_ _08817_ VPWR VGND _08820_ sg13g2_nor3_1
X_15935_ _08739_ _08818_ _08820_ VPWR VGND _08821_ sg13g2_a21o_1
X_15936_ _08739_ VPWR VGND _08822_ sg13g2_buf_1
X_15937_ _08822_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[17]\ VPWR VGND _08823_ sg13g2_nor2_1
X_15938_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2652_o\ _08821_ _08823_ _08817_ _08758_ VPWR 
+ VGND
+ _08824_ sg13g2_a221oi_1
X_15939_ _08762_ _07931_ _08824_ VPWR VGND _08825_ sg13g2_a21oi_1
X_15940_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2650_o[0]\ VPWR VGND _08826_ sg13g2_buf_1
X_15941_ _08826_ VPWR VGND _08827_ sg13g2_buf_1
X_15942_ _08825_ _08827_ VPWR VGND _08828_ sg13g2_nand2b_1
X_15943_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2652_o\ _08745_ VPWR VGND _08829_ sg13g2_nand2_1
X_15944_ _08740_ _08742_ _08829_ VPWR VGND _08830_ sg13g2_o21ai_1
X_15945_ _08830_ _08818_ VPWR VGND _08831_ sg13g2_nand2_1
X_15946_ _08819_ _08817_ VPWR VGND _08832_ sg13g2_and2_1
X_15947_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2652_o\ VPWR VGND _08833_ sg13g2_inv_1
X_15948_ _08819_ _08833_ _08817_ VPWR VGND _08834_ sg13g2_nor3_1
X_15949_ _08832_ _08834_ _08750_ VPWR VGND _08835_ sg13g2_o21ai_1
X_15950_ _08809_ _08813_ VPWR VGND _08836_ sg13g2_nor2_1
X_15951_ _08726_ _08763_ VPWR VGND _08837_ sg13g2_xor2_1
X_15952_ _08836_ _08837_ VPWR VGND _08838_ sg13g2_xnor2_1
X_15953_ _08729_ _08838_ VPWR VGND _08839_ sg13g2_nand2_1
X_15954_ _08651_ _08675_ VPWR VGND _08840_ sg13g2_xor2_1
X_15955_ _08840_ VPWR VGND _08841_ sg13g2_buf_1
X_15956_ _08795_ _08841_ VPWR VGND _08842_ sg13g2_xnor2_1
X_15957_ _08464_ VPWR VGND _08843_ sg13g2_buf_1
X_15958_ _08644_ VPWR VGND _08844_ sg13g2_buf_1
X_15959_ _08843_ _08844_ VPWR VGND _08845_ sg13g2_nand2_1
X_15960_ _08843_ _08845_ _08807_ VPWR VGND _08846_ sg13g2_mux2_1
X_15961_ _08793_ _08842_ _08846_ VPWR VGND _08847_ sg13g2_nand3_1
X_15962_ _08461_ VPWR VGND _08848_ sg13g2_inv_1
X_15963_ _08848_ VPWR VGND _08849_ sg13g2_buf_1
X_15964_ _08844_ _08807_ _08793_ VPWR VGND _08850_ sg13g2_o21ai_1
X_15965_ _08844_ _08793_ VPWR VGND _08851_ sg13g2_nor2_1
X_15966_ _08849_ _08850_ _08851_ VPWR VGND _08852_ sg13g2_a21oi_1
X_15967_ _08842_ _08852_ VPWR VGND _08853_ sg13g2_or2_1
X_15968_ _08568_ VPWR VGND _08854_ sg13g2_buf_1
X_15969_ _08781_ _08783_ _08785_ VPWR VGND _08855_ sg13g2_nor3_1
X_15970_ _08789_ _08855_ VPWR VGND _08856_ sg13g2_nor2_1
X_15971_ _08570_ _08766_ VPWR VGND _08857_ sg13g2_xnor2_1
X_15972_ _08856_ _08857_ VPWR VGND _08858_ sg13g2_xnor2_1
X_15973_ _08854_ _08858_ VPWR VGND _08859_ sg13g2_nand2_1
X_15974_ _08588_ VPWR VGND _08860_ sg13g2_inv_1
X_15975_ _08590_ VPWR VGND _08861_ sg13g2_buf_2
X_15976_ _08861_ _08778_ _08779_ VPWR VGND _08862_ sg13g2_a21oi_1
X_15977_ _08768_ _08862_ VPWR VGND _08863_ sg13g2_xor2_1
X_15978_ _08595_ _08863_ VPWR VGND _08864_ sg13g2_xnor2_1
X_15979_ _08860_ _08864_ VPWR VGND _08865_ sg13g2_nor2_1
X_15980_ _08635_ _08865_ VPWR VGND _08866_ sg13g2_nor2_1
X_15981_ _08578_ VPWR VGND _08867_ sg13g2_buf_2
X_15982_ _08867_ VPWR VGND _08868_ sg13g2_buf_1
X_15983_ _08868_ _08773_ _08774_ VPWR VGND _08869_ sg13g2_a21oi_1
X_15984_ _08551_ _08769_ VPWR VGND _08870_ sg13g2_xnor2_1
X_15985_ _08869_ _08870_ VPWR VGND _08871_ sg13g2_xnor2_1
X_15986_ _08527_ VPWR VGND _08872_ sg13g2_buf_1
X_15987_ _08542_ _08771_ VPWR VGND _08873_ sg13g2_nand2_1
X_15988_ _08867_ _08772_ VPWR VGND _08874_ sg13g2_xor2_1
X_15989_ _08873_ _08874_ VPWR VGND _08875_ sg13g2_xnor2_1
X_15990_ _08549_ _08871_ VPWR VGND _08876_ sg13g2_xor2_1
X_15991_ _08872_ _08875_ _08876_ VPWR VGND _08877_ sg13g2_a21oi_1
X_15992_ _08476_ VPWR VGND _08878_ sg13g2_buf_1
X_15993_ _08878_ VPWR VGND _08879_ sg13g2_buf_1
X_15994_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ VPWR VGND _08880_ sg13g2_inv_1
X_15995_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ VPWR VGND _08881_ sg13g2_inv_1
X_15996_ _08480_ VPWR VGND _08882_ sg13g2_buf_1
X_15997_ _08882_ VPWR VGND _08883_ sg13g2_buf_1
X_15998_ _08482_ VPWR VGND _08884_ sg13g2_buf_1
X_15999_ _08485_ VPWR VGND _08885_ sg13g2_buf_1
X_16000_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ VPWR VGND _08886_ sg13g2_inv_1
X_16001_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ VPWR VGND _08887_ sg13g2_inv_1
X_16002_ _08489_ VPWR VGND _08888_ sg13g2_buf_1
X_16003_ _08491_ VPWR VGND _08889_ sg13g2_buf_1
X_16004_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ VPWR VGND _08890_ sg13g2_buf_1
X_16005_ _08498_ VPWR VGND _08891_ sg13g2_buf_2
X_16006_ _08891_ VPWR VGND _08892_ sg13g2_buf_1
X_16007_ _08890_ _08892_ VPWR VGND _08893_ sg13g2_nand2b_1
X_16008_ _08494_ VPWR VGND _08894_ sg13g2_buf_1
X_16009_ _08894_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ VPWR VGND _08895_ sg13g2_nor2b_1
X_16010_ _08892_ _08890_ VPWR VGND _08896_ sg13g2_nor2b_1
X_16011_ _08889_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ _08893_ _08895_ _08896_ VPWR 
+ VGND
+ _08897_ sg13g2_a221oi_1
X_16012_ _08885_ _08886_ _08887_ _08888_ _08897_ VPWR 
+ VGND
+ _08898_ sg13g2_a221oi_1
X_16013_ _08487_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ _08884_ _08898_ VPWR 
+ VGND
+ _08899_ sg13g2_a221oi_1
X_16014_ _08879_ _08880_ _08881_ _08883_ _08899_ VPWR 
+ VGND
+ _08900_ sg13g2_a221oi_1
X_16015_ _08513_ _08473_ VPWR VGND _08901_ sg13g2_xnor2_1
X_16016_ _08771_ _08901_ VPWR VGND _08902_ sg13g2_xnor2_1
X_16017_ _08879_ _08880_ _08902_ VPWR VGND _08903_ sg13g2_o21ai_1
X_16018_ _08873_ _08874_ VPWR VGND _08904_ sg13g2_nor2_1
X_16019_ _08516_ _08874_ _08904_ VPWR VGND _08905_ sg13g2_a21oi_1
X_16020_ _08555_ VPWR VGND _08906_ sg13g2_inv_1
X_16021_ _08906_ VPWR VGND _08907_ sg13g2_buf_1
X_16022_ _08527_ _08907_ VPWR VGND _08908_ sg13g2_nand2_1
X_16023_ _08542_ _08771_ VPWR VGND _08909_ sg13g2_xnor2_1
X_16024_ _08908_ _08909_ VPWR VGND _08910_ sg13g2_nand2_1
X_16025_ _08872_ _08874_ _08910_ VPWR VGND _08911_ sg13g2_o21ai_1
X_16026_ _08557_ _08905_ _08911_ VPWR VGND _08912_ sg13g2_o21ai_1
X_16027_ _08900_ _08903_ _08912_ VPWR VGND _08913_ sg13g2_o21ai_1
X_16028_ _08605_ _08871_ _08877_ _08913_ VPWR VGND 
+ _08914_
+ sg13g2_a22oi_1
X_16029_ _08770_ _08776_ VPWR VGND _08915_ sg13g2_nor2_1
X_16030_ _08861_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[9]\ VPWR VGND _08916_ sg13g2_xnor2_1
X_16031_ _08915_ _08916_ VPWR VGND _08917_ sg13g2_xnor2_1
X_16032_ _08577_ _08917_ VPWR VGND _08918_ sg13g2_and2_1
X_16033_ _08574_ VPWR VGND _08919_ sg13g2_inv_1
X_16034_ _08919_ VPWR VGND _08920_ sg13g2_buf_1
X_16035_ _08920_ VPWR VGND _08921_ sg13g2_buf_1
X_16036_ _08917_ _08921_ VPWR VGND _08922_ sg13g2_nand2b_1
X_16037_ _08914_ _08918_ _08922_ VPWR VGND _08923_ sg13g2_o21ai_1
X_16038_ _08623_ _08863_ VPWR VGND _08924_ sg13g2_xor2_1
X_16039_ _08923_ _08924_ VPWR VGND _08925_ sg13g2_nand2_1
X_16040_ _08781_ _08783_ VPWR VGND _08926_ sg13g2_nor2_1
X_16041_ _08617_ _08784_ VPWR VGND _08927_ sg13g2_xnor2_1
X_16042_ _08926_ _08927_ VPWR VGND _08928_ sg13g2_xnor2_1
X_16043_ _08866_ _08925_ _08928_ VPWR VGND _08929_ sg13g2_a21oi_1
X_16044_ _08615_ VPWR VGND _08930_ sg13g2_buf_1
X_16045_ _08923_ _08924_ _08865_ VPWR VGND _08931_ sg13g2_a21oi_1
X_16046_ _08930_ _08931_ VPWR VGND _08932_ sg13g2_nor2_1
X_16047_ _08610_ _08858_ VPWR VGND _08933_ sg13g2_xnor2_1
X_16048_ _08929_ _08932_ _08933_ VPWR VGND _08934_ sg13g2_o21ai_1
X_16049_ _08847_ _08853_ _08859_ _08934_ VPWR VGND 
+ _08935_
+ sg13g2_a22oi_1
X_16050_ _08464_ _08811_ VPWR VGND _08936_ sg13g2_and2_1
X_16051_ _08811_ _08807_ _08936_ _08793_ VPWR VGND 
+ _08937_
+ sg13g2_a22oi_1
X_16052_ _08937_ VPWR VGND _08938_ sg13g2_buf_1
X_16053_ _08796_ _08938_ VPWR VGND _08939_ sg13g2_nand2_1
X_16054_ _08668_ VPWR VGND _08940_ sg13g2_buf_1
X_16055_ _08940_ _08794_ VPWR VGND _08941_ sg13g2_xor2_1
X_16056_ _08939_ _08941_ VPWR VGND _08942_ sg13g2_xor2_1
X_16057_ _08684_ VPWR VGND _08943_ sg13g2_buf_1
X_16058_ _08843_ _08793_ VPWR VGND _08944_ sg13g2_and2_1
X_16059_ _08944_ _08807_ VPWR VGND _08945_ sg13g2_nor2_1
X_16060_ _08811_ _08796_ VPWR VGND _08946_ sg13g2_nand2_1
X_16061_ _08945_ _08946_ VPWR VGND _08947_ sg13g2_xnor2_1
X_16062_ _08793_ _08842_ VPWR VGND _08948_ sg13g2_nor2_1
X_16063_ _08807_ _08842_ _08948_ VPWR VGND _08949_ sg13g2_a21oi_1
X_16064_ _08807_ _08842_ _08944_ VPWR VGND _08950_ sg13g2_nand3b_1
X_16065_ _08843_ _08949_ _08950_ VPWR VGND _08951_ sg13g2_o21ai_1
X_16066_ _08943_ _08947_ _08951_ _08646_ VPWR VGND 
+ _08952_
+ sg13g2_a22oi_1
X_16067_ _08681_ _08942_ _08952_ VPWR VGND _08953_ sg13g2_o21ai_1
X_16068_ _08679_ VPWR VGND _08954_ sg13g2_inv_1
X_16069_ _08954_ VPWR VGND _08955_ sg13g2_buf_1
X_16070_ _08794_ _08939_ VPWR VGND _08956_ sg13g2_nor2_1
X_16071_ _08682_ _08795_ VPWR VGND _08957_ sg13g2_and2_1
X_16072_ _08940_ _08794_ _08957_ VPWR VGND _08958_ sg13g2_nor3_1
X_16073_ _08955_ _08956_ _08958_ _08938_ VPWR VGND 
+ _08959_
+ sg13g2_a22oi_1
X_16074_ _08696_ _08954_ VPWR VGND _08960_ sg13g2_nand2_1
X_16075_ _08957_ _08960_ VPWR VGND _08961_ sg13g2_nor2_1
X_16076_ _08763_ _08704_ VPWR VGND _08962_ sg13g2_xnor2_1
X_16077_ _08794_ _08960_ _08962_ VPWR VGND _08963_ sg13g2_o21ai_1
X_16078_ _08938_ _08961_ _08963_ VPWR VGND _08964_ sg13g2_a21oi_1
X_16079_ _08940_ _08794_ VPWR VGND _08965_ sg13g2_and2_1
X_16080_ _08680_ _08939_ VPWR VGND _08966_ sg13g2_nand2_1
X_16081_ _08939_ _08941_ _08965_ _08966_ _08962_ VPWR 
+ VGND
+ _08967_ sg13g2_a221oi_1
X_16082_ _08959_ _08964_ _08967_ VPWR VGND _08968_ sg13g2_a21oi_1
X_16083_ _08935_ _08953_ _08968_ VPWR VGND _08969_ sg13g2_o21ai_1
X_16084_ _08758_ VPWR VGND _08970_ sg13g2_buf_1
X_16085_ _08831_ _08835_ _08839_ _08969_ _08970_ VPWR 
+ VGND
+ _08971_ sg13g2_a221oi_1
X_16086_ _08761_ _08828_ _08971_ VPWR VGND _00494_ sg13g2_a21oi_1
X_16087_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2650_o[1]\ VPWR VGND _08972_ sg13g2_buf_1
X_16088_ _08972_ VPWR VGND _08973_ sg13g2_inv_1
X_16089_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2647_o[1]\ VPWR VGND _08974_ sg13g2_buf_1
X_16090_ _08974_ _08759_ VPWR VGND _08975_ sg13g2_nand2_1
X_16091_ _08973_ _08825_ _08975_ VPWR VGND _08976_ sg13g2_o21ai_1
X_16092_ _08971_ _08976_ VPWR VGND _00495_ sg13g2_nor2b_1
X_16093_ _07931_ VPWR VGND _08977_ sg13g2_buf_1
X_16094_ _08827_ _08977_ VPWR VGND _08978_ sg13g2_nor2_1
X_16095_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2653_o[0]\ VPWR VGND _08979_ sg13g2_buf_2
X_16096_ _08979_ VPWR VGND _08980_ sg13g2_buf_2
X_16097_ _08759_ VPWR VGND _08981_ sg13g2_buf_1
X_16098_ _08980_ _08981_ VPWR VGND _08982_ sg13g2_nor2_1
X_16099_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[16]\ VPWR VGND _08983_ sg13g2_buf_1
X_16100_ _08983_ VPWR VGND _08984_ sg13g2_inv_1
X_16101_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[15]\ VPWR VGND _08985_ sg13g2_buf_1
X_16102_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[13]\ VPWR VGND _08986_ sg13g2_buf_1
X_16103_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[11]\ VPWR VGND _08987_ sg13g2_buf_1
X_16104_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[12]\ VPWR VGND _08988_ sg13g2_buf_1
X_16105_ _08454_ _08988_ VPWR VGND _08989_ sg13g2_nand2_1
X_16106_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[10]\ VPWR VGND _08990_ sg13g2_buf_1
X_16107_ _08594_ _08990_ VPWR VGND _08991_ sg13g2_nand2_1
X_16108_ _08989_ _08991_ VPWR VGND _08992_ sg13g2_nand2_1
X_16109_ _08987_ _08992_ VPWR VGND _08993_ sg13g2_nor2_1
X_16110_ _08406_ VPWR VGND _08994_ sg13g2_buf_1
X_16111_ _08994_ _08992_ VPWR VGND _08995_ sg13g2_nor2_1
X_16112_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[9]\ VPWR VGND _08996_ sg13g2_buf_1
X_16113_ _08996_ VPWR VGND _08997_ sg13g2_inv_1
X_16114_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[8]\ VPWR VGND _08998_ sg13g2_buf_1
X_16115_ _08436_ _08998_ VPWR VGND _08999_ sg13g2_nor2_1
X_16116_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[6]\ VPWR VGND _09000_ sg13g2_buf_1
X_16117_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[7]\ VPWR VGND _09001_ sg13g2_buf_1
X_16118_ _08426_ _09000_ _09001_ VPWR VGND _09002_ sg13g2_a21o_1
X_16119_ _08426_ _09001_ _09000_ VPWR VGND _09003_ sg13g2_and3_1
X_16120_ _08417_ _08998_ _09002_ _08422_ _09003_ VPWR 
+ VGND
+ _09004_ sg13g2_a221oi_1
X_16121_ _09004_ VPWR VGND _09005_ sg13g2_buf_1
X_16122_ _08997_ _08999_ _09005_ VPWR VGND _09006_ sg13g2_nor3_1
X_16123_ _08999_ _09005_ _08997_ VPWR VGND _09007_ sg13g2_o21ai_1
X_16124_ _08413_ _09006_ _09007_ VPWR VGND _09008_ sg13g2_o21ai_1
X_16125_ _09008_ VPWR VGND _09009_ sg13g2_buf_1
X_16126_ _08993_ _08995_ _09009_ VPWR VGND _09010_ sg13g2_o21ai_1
X_16127_ _08994_ _08987_ VPWR VGND _09011_ sg13g2_nor2_1
X_16128_ _08594_ _08990_ VPWR VGND _09012_ sg13g2_nor2_1
X_16129_ _08989_ _09012_ VPWR VGND _09013_ sg13g2_nand2_1
X_16130_ _08408_ _08987_ _09013_ VPWR VGND _09014_ sg13g2_a21oi_1
X_16131_ _08989_ _09011_ _09014_ VPWR VGND _09015_ sg13g2_a21oi_1
X_16132_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[14]\ VPWR VGND _09016_ sg13g2_buf_1
X_16133_ _08651_ _09016_ VPWR VGND _09017_ sg13g2_nor2_1
X_16134_ _08455_ _08988_ VPWR VGND _09018_ sg13g2_or2_1
X_16135_ _09017_ _09018_ VPWR VGND _09019_ sg13g2_nor2b_1
X_16136_ _08986_ _09010_ _09015_ _09019_ VPWR VGND 
+ _09020_
+ sg13g2_nand4_1
X_16137_ _08463_ _09010_ _09015_ _09019_ VPWR VGND 
+ _09021_
+ sg13g2_nand4_1
X_16138_ _08462_ _08986_ VPWR VGND _09022_ sg13g2_nand2_1
X_16139_ _09017_ _09022_ VPWR VGND _09023_ sg13g2_nor2_1
X_16140_ _08652_ _09016_ _09023_ VPWR VGND _09024_ sg13g2_a21oi_1
X_16141_ _09020_ _09021_ _09024_ VPWR VGND _09025_ sg13g2_nand3_1
X_16142_ _09025_ VPWR VGND _09026_ sg13g2_buf_1
X_16143_ _08985_ _09026_ VPWR VGND _09027_ sg13g2_nand2_1
X_16144_ _08985_ _09026_ _08668_ VPWR VGND _09028_ sg13g2_o21ai_1
X_16145_ _08716_ _08984_ _09027_ _09028_ VPWR VGND 
+ _09029_
+ sg13g2_a22oi_1
X_16146_ _08726_ _08983_ _09029_ VPWR VGND _09030_ sg13g2_a21oi_1
X_16147_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[17]\ VPWR VGND _09031_ sg13g2_buf_1
X_16148_ _08738_ _09031_ VPWR VGND _09032_ sg13g2_xor2_1
X_16149_ _09030_ _09032_ VPWR VGND _09033_ sg13g2_xnor2_1
X_16150_ _08744_ _09033_ VPWR VGND _09034_ sg13g2_xnor2_1
X_16151_ _08728_ VPWR VGND _09035_ sg13g2_inv_1
X_16152_ _09027_ _09028_ VPWR VGND _09036_ sg13g2_nand2_1
X_16153_ _08983_ _09036_ VPWR VGND _09037_ sg13g2_xnor2_1
X_16154_ _08726_ _09037_ VPWR VGND _09038_ sg13g2_xnor2_1
X_16155_ _09035_ _09038_ VPWR VGND _09039_ sg13g2_nor2_1
X_16156_ _08762_ _09033_ VPWR VGND _09040_ sg13g2_nor2_1
X_16157_ _09034_ _09039_ _09040_ VPWR VGND _09041_ sg13g2_a21oi_1
X_16158_ _09009_ _08991_ _09012_ VPWR VGND _09042_ sg13g2_a21oi_1
X_16159_ _08616_ _08987_ VPWR VGND _09043_ sg13g2_or2_1
X_16160_ _08616_ _08987_ VPWR VGND _09044_ sg13g2_and2_1
X_16161_ _09042_ _09043_ _09044_ VPWR VGND _09045_ sg13g2_a21oi_1
X_16162_ _08570_ _08988_ VPWR VGND _09046_ sg13g2_xnor2_1
X_16163_ _09045_ _09046_ VPWR VGND _09047_ sg13g2_xnor2_1
X_16164_ _08589_ VPWR VGND _09048_ sg13g2_buf_1
X_16165_ _08595_ _08990_ VPWR VGND _09049_ sg13g2_xnor2_1
X_16166_ _09009_ _09049_ VPWR VGND _09050_ sg13g2_xnor2_1
X_16167_ _09048_ _09050_ _08635_ VPWR VGND _09051_ sg13g2_a21oi_1
X_16168_ _09048_ _09050_ VPWR VGND _09052_ sg13g2_nand2_1
X_16169_ _08617_ _08987_ VPWR VGND _09053_ sg13g2_xnor2_1
X_16170_ _09042_ _09053_ VPWR VGND _09054_ sg13g2_xnor2_1
X_16171_ _09052_ _09054_ VPWR VGND _09055_ sg13g2_and2_1
X_16172_ _08543_ _09000_ VPWR VGND _09056_ sg13g2_nand2_1
X_16173_ _08868_ _09001_ VPWR VGND _09057_ sg13g2_xor2_1
X_16174_ _09056_ _09057_ VPWR VGND _09058_ sg13g2_xnor2_1
X_16175_ _08514_ _09000_ VPWR VGND _09059_ sg13g2_xnor2_1
X_16176_ _08474_ _09059_ VPWR VGND _09060_ sg13g2_xnor2_1
X_16177_ _08477_ VPWR VGND _09061_ sg13g2_buf_1
X_16178_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[119]\ VPWR VGND _09062_ sg13g2_buf_1
X_16179_ _09061_ _09062_ VPWR VGND _09063_ sg13g2_nor2_1
X_16180_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ VPWR VGND _09064_ sg13g2_buf_1
X_16181_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ VPWR VGND _09065_ sg13g2_buf_1
X_16182_ _08482_ _09065_ VPWR VGND _09066_ sg13g2_nand2_1
X_16183_ _09064_ _09066_ VPWR VGND _09067_ sg13g2_nand2b_1
X_16184_ _08485_ _09066_ VPWR VGND _09068_ sg13g2_nand2_1
X_16185_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ VPWR VGND _09069_ sg13g2_inv_1
X_16186_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[115]\ VPWR VGND _09070_ sg13g2_buf_1
X_16187_ _08498_ VPWR VGND _09071_ sg13g2_buf_1
X_16188_ _09070_ _09071_ VPWR VGND _09072_ sg13g2_nand2b_1
X_16189_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ VPWR VGND _09073_ sg13g2_nor2b_1
X_16190_ _09071_ _09070_ VPWR VGND _09074_ sg13g2_nor2b_1
X_16191_ _08491_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _09072_ _09073_ _09074_ VPWR 
+ VGND
+ _09075_ sg13g2_a221oi_1
X_16192_ _08888_ _09069_ _09075_ VPWR VGND _09076_ sg13g2_a21oi_1
X_16193_ _09067_ _09068_ _09076_ VPWR VGND _09077_ sg13g2_a21o_1
X_16194_ _08487_ _09064_ VPWR VGND _09078_ sg13g2_nor2_1
X_16195_ _08482_ _09065_ VPWR VGND _09079_ sg13g2_nor2_1
X_16196_ _09066_ _09078_ _09079_ VPWR VGND _09080_ sg13g2_a21oi_1
X_16197_ _09062_ _09060_ VPWR VGND _09081_ sg13g2_nand2b_1
X_16198_ _08878_ _09060_ VPWR VGND _09082_ sg13g2_nand2_1
X_16199_ _09077_ _09080_ _09081_ _09082_ VPWR VGND 
+ _09083_
+ sg13g2_a22oi_1
X_16200_ _08557_ _09059_ _09060_ _09063_ _09083_ VPWR 
+ VGND
+ _09084_ sg13g2_a221oi_1
X_16201_ _09058_ _09084_ _08872_ VPWR VGND _09085_ sg13g2_a21oi_1
X_16202_ _08868_ _09002_ _09003_ VPWR VGND _09086_ sg13g2_a21oi_1
X_16203_ _08551_ _08998_ VPWR VGND _09087_ sg13g2_xnor2_1
X_16204_ _09086_ _09087_ VPWR VGND _09088_ sg13g2_xnor2_1
X_16205_ _08999_ _09005_ VPWR VGND _09089_ sg13g2_nor2_1
X_16206_ _08584_ _08996_ VPWR VGND _09090_ sg13g2_xor2_1
X_16207_ _09089_ _09090_ VPWR VGND _09091_ sg13g2_xnor2_1
X_16208_ _08605_ _09088_ _09091_ _08921_ VPWR VGND 
+ _09092_
+ sg13g2_a22oi_1
X_16209_ _09058_ _09084_ _09092_ VPWR VGND _09093_ sg13g2_o21ai_1
X_16210_ _08861_ _08996_ VPWR VGND _09094_ sg13g2_nand2_1
X_16211_ _08577_ _09089_ _09094_ VPWR VGND _09095_ sg13g2_a21oi_1
X_16212_ _09089_ _09090_ _09095_ VPWR VGND _09096_ sg13g2_a21oi_1
X_16213_ _08990_ _08623_ VPWR VGND _09097_ sg13g2_xor2_1
X_16214_ _08549_ _09088_ VPWR VGND _09098_ sg13g2_xor2_1
X_16215_ _08996_ _09089_ VPWR VGND _09099_ sg13g2_nor2_1
X_16216_ _08577_ _09006_ _09007_ VPWR VGND _09100_ sg13g2_o21ai_1
X_16217_ _08921_ _09099_ _09100_ _08625_ _09097_ VPWR 
+ VGND
+ _09101_ sg13g2_a221oi_1
X_16218_ _09096_ _09097_ _09092_ _09098_ _09101_ VPWR 
+ VGND
+ _09102_ sg13g2_a221oi_1
X_16219_ _09085_ _09093_ _09102_ VPWR VGND _09103_ sg13g2_o21ai_1
X_16220_ _09051_ _09055_ _09103_ VPWR VGND _09104_ sg13g2_o21ai_1
X_16221_ _08610_ VPWR VGND _09105_ sg13g2_inv_1
X_16222_ _09105_ VPWR VGND _09106_ sg13g2_buf_1
X_16223_ _09106_ _09047_ VPWR VGND _09107_ sg13g2_xnor2_1
X_16224_ _08930_ _09054_ _09107_ VPWR VGND _09108_ sg13g2_a21oi_1
X_16225_ _09010_ _09015_ _09018_ VPWR VGND _09109_ sg13g2_and3_1
X_16226_ _09109_ VPWR VGND _09110_ sg13g2_buf_1
X_16227_ _08464_ _08986_ VPWR VGND _09111_ sg13g2_xor2_1
X_16228_ _09110_ _09111_ VPWR VGND _09112_ sg13g2_xor2_1
X_16229_ _08844_ _09112_ VPWR VGND _09113_ sg13g2_nor2_1
X_16230_ _08854_ _09047_ _09104_ _09108_ _09113_ VPWR 
+ VGND
+ _09114_ sg13g2_a221oi_1
X_16231_ _08986_ _09110_ VPWR VGND _09115_ sg13g2_nor2_1
X_16232_ _08986_ _09110_ VPWR VGND _09116_ sg13g2_nand2_1
X_16233_ _08645_ _09116_ _09115_ VPWR VGND _09117_ sg13g2_a21o_1
X_16234_ _08646_ _09115_ _09117_ _08849_ VPWR VGND 
+ _09118_
+ sg13g2_a22oi_1
X_16235_ _08644_ _09110_ _09022_ VPWR VGND _09119_ sg13g2_a21oi_1
X_16236_ _09110_ _09111_ _09119_ VPWR VGND _09120_ sg13g2_a21oi_1
X_16237_ _09016_ _08841_ VPWR VGND _09121_ sg13g2_xnor2_1
X_16238_ _09118_ _09120_ _09121_ VPWR VGND _09122_ sg13g2_mux2_1
X_16239_ _09114_ _09122_ VPWR VGND _09123_ sg13g2_or2_1
X_16240_ _08849_ _09116_ _09115_ VPWR VGND _09124_ sg13g2_a21oi_1
X_16241_ _08682_ _09016_ VPWR VGND _09125_ sg13g2_xor2_1
X_16242_ _09124_ _09125_ VPWR VGND _09126_ sg13g2_xnor2_1
X_16243_ _08940_ _08985_ VPWR VGND _09127_ sg13g2_xor2_1
X_16244_ _09026_ _09127_ VPWR VGND _09128_ sg13g2_xnor2_1
X_16245_ _08943_ _09126_ _09128_ VPWR VGND _09129_ sg13g2_a21oi_1
X_16246_ _09123_ _09129_ _08681_ VPWR VGND _09130_ sg13g2_a21oi_1
X_16247_ _08684_ _09126_ VPWR VGND _09131_ sg13g2_nand2_1
X_16248_ _09114_ _09122_ _09131_ VPWR VGND _09132_ sg13g2_o21ai_1
X_16249_ _09128_ _09132_ VPWR VGND _09133_ sg13g2_and2_1
X_16250_ _09031_ _08750_ VPWR VGND _09134_ sg13g2_xnor2_1
X_16251_ _08983_ _09036_ _09134_ VPWR VGND _09135_ sg13g2_nor3_1
X_16252_ _08983_ _09036_ _09134_ VPWR VGND _09136_ sg13g2_nand3_1
X_16253_ _09135_ _09136_ VPWR VGND _09137_ sg13g2_nor2b_1
X_16254_ _08726_ _08702_ _09134_ VPWR VGND _09138_ sg13g2_nand3_1
X_16255_ _08726_ _08702_ _09134_ VPWR VGND _09139_ sg13g2_or3_1
X_16256_ _09138_ _09139_ _09037_ VPWR VGND _09140_ sg13g2_a21o_1
X_16257_ _08704_ _09137_ _09140_ VPWR VGND _09141_ sg13g2_o21ai_1
X_16258_ _09130_ _09133_ _09141_ VPWR VGND _09142_ sg13g2_o21ai_1
X_16259_ _09031_ VPWR VGND _09143_ sg13g2_inv_1
X_16260_ _09143_ _09030_ _08712_ VPWR VGND _09144_ sg13g2_a21oi_1
X_16261_ _09143_ _09030_ VPWR VGND _09145_ sg13g2_nor2_1
X_16262_ _09144_ _09145_ VPWR VGND _09146_ sg13g2_nor2_1
X_16263_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2655_o\ _09146_ _07931_ VPWR VGND _09147_ sg13g2_o21ai_1
X_16264_ _09041_ _09142_ _09147_ VPWR VGND _09148_ sg13g2_a21oi_1
X_16265_ _08978_ _08982_ _09148_ VPWR VGND _00496_ sg13g2_nor3_1
X_16266_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2653_o[1]\ VPWR VGND _09149_ sg13g2_buf_2
X_16267_ _09149_ VPWR VGND _09150_ sg13g2_buf_2
X_16268_ _07931_ VPWR VGND _09151_ sg13g2_buf_1
X_16269_ _08973_ _07932_ VPWR VGND _09152_ sg13g2_nor2_1
X_16270_ _09150_ _09151_ _09152_ VPWR VGND _09153_ sg13g2_a21oi_1
X_16271_ _09148_ _09153_ VPWR VGND _00497_ sg13g2_nor2_1
X_16272_ _08970_ VPWR VGND _09154_ sg13g2_buf_1
X_16273_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[17]\ VPWR VGND _09155_ sg13g2_buf_1
X_16274_ _08710_ _09155_ VPWR VGND _09156_ sg13g2_nor2_1
X_16275_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2658_o\ VPWR VGND _09157_ sg13g2_buf_1
X_16276_ _08822_ _09155_ _09157_ VPWR VGND _09158_ sg13g2_and3_1
X_16277_ _08741_ _07801_ VPWR VGND _09159_ sg13g2_nand2_1
X_16278_ _09157_ _09156_ _08707_ VPWR VGND _09160_ sg13g2_o21ai_1
X_16279_ _08744_ _07801_ _09160_ VPWR VGND _09161_ sg13g2_nand3_1
X_16280_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[16]\ VPWR VGND _09162_ sg13g2_buf_1
X_16281_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[15]\ VPWR VGND _09163_ sg13g2_buf_1
X_16282_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[13]\ VPWR VGND _09164_ sg13g2_buf_1
X_16283_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[11]\ VPWR VGND _09165_ sg13g2_buf_1
X_16284_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[12]\ VPWR VGND _09166_ sg13g2_buf_1
X_16285_ _08453_ _09166_ VPWR VGND _09167_ sg13g2_nor2_1
X_16286_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[10]\ VPWR VGND _09168_ sg13g2_buf_1
X_16287_ _08594_ _09168_ VPWR VGND _09169_ sg13g2_nor2_1
X_16288_ _09167_ _09169_ VPWR VGND _09170_ sg13g2_nor2_1
X_16289_ _09165_ _09170_ VPWR VGND _09171_ sg13g2_nand2_1
X_16290_ _08994_ _09170_ VPWR VGND _09172_ sg13g2_nand2_1
X_16291_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[8]\ VPWR VGND _09173_ sg13g2_buf_1
X_16292_ _08436_ _09173_ VPWR VGND _09174_ sg13g2_nor2_1
X_16293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[6]\ VPWR VGND _09175_ sg13g2_buf_1
X_16294_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[7]\ VPWR VGND _09176_ sg13g2_buf_1
X_16295_ _08426_ _09175_ _09176_ VPWR VGND _09177_ sg13g2_a21o_1
X_16296_ _08426_ _09176_ _09175_ VPWR VGND _09178_ sg13g2_and3_1
X_16297_ _08417_ _09173_ _09177_ _08422_ _09178_ VPWR 
+ VGND
+ _09179_ sg13g2_a221oi_1
X_16298_ _09179_ VPWR VGND _09180_ sg13g2_buf_1
X_16299_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[9]\ VPWR VGND _09181_ sg13g2_buf_1
X_16300_ _09181_ VPWR VGND _09182_ sg13g2_inv_1
X_16301_ _09174_ _09180_ _09182_ VPWR VGND _09183_ sg13g2_o21ai_1
X_16302_ _09182_ _09174_ _09180_ VPWR VGND _09184_ sg13g2_nor3_1
X_16303_ _08582_ _09183_ _09184_ VPWR VGND _09185_ sg13g2_a21oi_1
X_16304_ _09171_ _09172_ _09185_ VPWR VGND _09186_ sg13g2_a21oi_1
X_16305_ _08407_ _09165_ VPWR VGND _09187_ sg13g2_nand2_1
X_16306_ _08594_ _09168_ VPWR VGND _09188_ sg13g2_nand2_1
X_16307_ _09167_ _09188_ VPWR VGND _09189_ sg13g2_nor2_1
X_16308_ _08407_ _09165_ _09189_ VPWR VGND _09190_ sg13g2_o21ai_1
X_16309_ _09167_ _09187_ _09190_ VPWR VGND _09191_ sg13g2_o21ai_1
X_16310_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[14]\ VPWR VGND _09192_ sg13g2_buf_1
X_16311_ _08651_ _09192_ VPWR VGND _09193_ sg13g2_nand2_1
X_16312_ _08455_ _09166_ VPWR VGND _09194_ sg13g2_nand2_1
X_16313_ _09193_ _09194_ VPWR VGND _09195_ sg13g2_nand2_1
X_16314_ _09164_ _09186_ _09191_ _09195_ VPWR VGND 
+ _09196_
+ sg13g2_nor4_1
X_16315_ _08462_ _09186_ _09191_ _09195_ VPWR VGND 
+ _09197_
+ sg13g2_nor4_1
X_16316_ _09164_ VPWR VGND _09198_ sg13g2_inv_1
X_16317_ _08848_ _09198_ _09193_ VPWR VGND _09199_ sg13g2_nand3_1
X_16318_ _08652_ _09192_ _09199_ VPWR VGND _09200_ sg13g2_o21ai_1
X_16319_ _09196_ _09197_ _09200_ VPWR VGND _09201_ sg13g2_nor3_1
X_16320_ _09201_ VPWR VGND _09202_ sg13g2_buf_1
X_16321_ _09163_ _09202_ VPWR VGND _09203_ sg13g2_nor2_1
X_16322_ _09163_ _09202_ _08668_ VPWR VGND _09204_ sg13g2_a21oi_1
X_16323_ _08701_ VPWR VGND _09205_ sg13g2_buf_1
X_16324_ _09205_ _09162_ VPWR VGND _09206_ sg13g2_nand2_1
X_16325_ _09203_ _09204_ _09206_ VPWR VGND _09207_ sg13g2_o21ai_1
X_16326_ _08725_ _09162_ _09207_ VPWR VGND _09208_ sg13g2_o21ai_1
X_16327_ _09208_ VPWR VGND _09209_ sg13g2_buf_1
X_16328_ _09159_ _09161_ _09209_ VPWR VGND _09210_ sg13g2_mux2_1
X_16329_ _09156_ _09158_ _09210_ VPWR VGND _09211_ sg13g2_o21ai_1
X_16330_ _08738_ _09155_ VPWR VGND _09212_ sg13g2_xor2_1
X_16331_ _09157_ _09161_ VPWR VGND _09213_ sg13g2_and2_1
X_16332_ _09213_ _09159_ _09209_ VPWR VGND _09214_ sg13g2_mux2_1
X_16333_ _09161_ _09159_ _09212_ _09214_ VPWR VGND 
+ _09215_
+ sg13g2_a22oi_1
X_16334_ _09211_ _09215_ VPWR VGND _09216_ sg13g2_nand2_1
X_16335_ _09212_ _09209_ VPWR VGND _09217_ sg13g2_xnor2_1
X_16336_ _09217_ _08708_ VPWR VGND _09218_ sg13g2_nand2b_1
X_16337_ _08669_ _09163_ VPWR VGND _09219_ sg13g2_xor2_1
X_16338_ _09202_ _09219_ VPWR VGND _09220_ sg13g2_xnor2_1
X_16339_ _09191_ VPWR VGND _09221_ sg13g2_inv_1
X_16340_ _09186_ _09221_ _09194_ VPWR VGND _09222_ sg13g2_nand3b_1
X_16341_ _09222_ VPWR VGND _09223_ sg13g2_buf_1
X_16342_ _09164_ _09223_ _08464_ VPWR VGND _09224_ sg13g2_a21o_1
X_16343_ _09164_ _09223_ _09224_ VPWR VGND _09225_ sg13g2_o21ai_1
X_16344_ _09192_ _09225_ VPWR VGND _09226_ sg13g2_xor2_1
X_16345_ _08686_ _09226_ VPWR VGND _09227_ sg13g2_xnor2_1
X_16346_ _08955_ _09220_ _09227_ _08943_ VPWR VGND 
+ _09228_
+ sg13g2_a22oi_1
X_16347_ _08844_ VPWR VGND _09229_ sg13g2_buf_1
X_16348_ _09185_ _09169_ _09188_ VPWR VGND _09230_ sg13g2_o21ai_1
X_16349_ _09230_ VPWR VGND _09231_ sg13g2_buf_1
X_16350_ _08408_ _09165_ VPWR VGND _09232_ sg13g2_xnor2_1
X_16351_ _09231_ _09232_ VPWR VGND _09233_ sg13g2_xnor2_1
X_16352_ _08595_ _09168_ VPWR VGND _09234_ sg13g2_xnor2_1
X_16353_ _09185_ _09234_ VPWR VGND _09235_ sg13g2_xnor2_1
X_16354_ _08589_ _09235_ VPWR VGND _09236_ sg13g2_nand2_1
X_16355_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[138]\ VPWR VGND _09237_ sg13g2_buf_1
X_16356_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ VPWR VGND _09238_ sg13g2_inv_1
X_16357_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ VPWR VGND _09239_ sg13g2_inv_1
X_16358_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ VPWR VGND _09240_ sg13g2_buf_1
X_16359_ _09240_ _08489_ VPWR VGND _09241_ sg13g2_nand2b_1
X_16360_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ VPWR VGND _09242_ sg13g2_buf_1
X_16361_ _09242_ _08498_ VPWR VGND _09243_ sg13g2_nor2b_1
X_16362_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ VPWR VGND _09244_ sg13g2_nand2b_1
X_16363_ _08891_ _09242_ VPWR VGND _09245_ sg13g2_nand2b_1
X_16364_ _09243_ _09244_ _09245_ VPWR VGND _09246_ sg13g2_o21ai_1
X_16365_ _08888_ _09240_ VPWR VGND _09247_ sg13g2_nor2b_1
X_16366_ _08486_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ _09241_ _09246_ _09247_ VPWR 
+ VGND
+ _09248_ sg13g2_a221oi_1
X_16367_ _08885_ _09238_ _09239_ _08883_ _09248_ VPWR 
+ VGND
+ _09249_ sg13g2_a221oi_1
X_16368_ _09061_ _09237_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ _08482_ _09249_ VPWR 
+ VGND
+ _09250_ sg13g2_a221oi_1
X_16369_ _08469_ _09176_ VPWR VGND _09251_ sg13g2_xor2_1
X_16370_ _09251_ VPWR VGND _09252_ sg13g2_buf_1
X_16371_ _08527_ _09252_ VPWR VGND _09253_ sg13g2_nor2_1
X_16372_ _08542_ _09175_ VPWR VGND _09254_ sg13g2_xnor2_1
X_16373_ _09253_ _09254_ _08908_ VPWR VGND _09255_ sg13g2_o21ai_1
X_16374_ _09175_ VPWR VGND _09256_ sg13g2_inv_1
X_16375_ _08515_ _09256_ _09252_ VPWR VGND _09257_ sg13g2_nor3_1
X_16376_ _08515_ _09252_ _09257_ VPWR VGND _09258_ sg13g2_a21oi_1
X_16377_ _08556_ _09258_ VPWR VGND _09259_ sg13g2_nor2_1
X_16378_ _09237_ _08878_ VPWR VGND _09260_ sg13g2_nand2b_1
X_16379_ _09255_ _09259_ _09260_ VPWR VGND _09261_ sg13g2_o21ai_1
X_16380_ _08578_ _09177_ _09178_ VPWR VGND _09262_ sg13g2_a21oi_1
X_16381_ _08550_ _09173_ VPWR VGND _09263_ sg13g2_xnor2_1
X_16382_ _09262_ _09263_ VPWR VGND _09264_ sg13g2_xnor2_1
X_16383_ _08548_ _09264_ VPWR VGND _09265_ sg13g2_xor2_1
X_16384_ _08527_ _09252_ VPWR VGND _09266_ sg13g2_nand2_1
X_16385_ _09175_ _09266_ VPWR VGND _09267_ sg13g2_nor2_1
X_16386_ _09253_ _08474_ _09256_ VPWR VGND _09268_ sg13g2_nand3b_1
X_16387_ _08473_ _08555_ VPWR VGND _09269_ sg13g2_or2_1
X_16388_ _09269_ VPWR VGND _09270_ sg13g2_buf_1
X_16389_ _09252_ _09270_ _08532_ VPWR VGND _09271_ sg13g2_a21oi_1
X_16390_ _09252_ _09270_ VPWR VGND _09272_ sg13g2_nor2_1
X_16391_ _09271_ _09272_ _09175_ VPWR VGND _09273_ sg13g2_o21ai_1
X_16392_ _09268_ _09273_ _08516_ VPWR VGND _09274_ sg13g2_a21oi_1
X_16393_ _08473_ _08555_ _09175_ VPWR VGND _09275_ sg13g2_nor3_1
X_16394_ _08474_ _09175_ _09275_ VPWR VGND _09276_ sg13g2_a21oi_1
X_16395_ _09253_ _09276_ _09266_ VPWR VGND _09277_ sg13g2_o21ai_1
X_16396_ _08516_ _09277_ VPWR VGND _09278_ sg13g2_and2_1
X_16397_ _09265_ _09267_ _09274_ _09278_ VPWR VGND 
+ _09279_
+ sg13g2_nor4_1
X_16398_ _09250_ _09261_ _09279_ VPWR VGND _09280_ sg13g2_o21ai_1
X_16399_ _09174_ _09180_ VPWR VGND _09281_ sg13g2_nor2_1
X_16400_ _08583_ _09181_ VPWR VGND _09282_ sg13g2_xor2_1
X_16401_ _09281_ _09282_ VPWR VGND _09283_ sg13g2_xnor2_1
X_16402_ _08605_ _09264_ _09283_ _08921_ VPWR VGND 
+ _09284_
+ sg13g2_a22oi_1
X_16403_ _09233_ _09236_ _09280_ _09284_ VPWR VGND 
+ _09285_
+ sg13g2_nand4_1
X_16404_ _08615_ _09236_ _09280_ _09284_ VPWR VGND 
+ _09286_
+ sg13g2_nand4_1
X_16405_ _08584_ _09181_ VPWR VGND _09287_ sg13g2_nand2_1
X_16406_ _08576_ _09281_ _09287_ VPWR VGND _09288_ sg13g2_a21oi_1
X_16407_ _09281_ _09282_ _09288_ VPWR VGND _09289_ sg13g2_a21oi_1
X_16408_ _09168_ _08623_ VPWR VGND _09290_ sg13g2_xor2_1
X_16409_ _09181_ _09281_ VPWR VGND _09291_ sg13g2_nor2_1
X_16410_ _08576_ _09184_ _09183_ VPWR VGND _09292_ sg13g2_o21ai_1
X_16411_ _08920_ _09291_ _09292_ _08625_ _09290_ VPWR 
+ VGND
+ _09293_ sg13g2_a221oi_1
X_16412_ _09289_ _09290_ _09293_ VPWR VGND _09294_ sg13g2_a21o_1
X_16413_ _09233_ _09236_ _09294_ VPWR VGND _09295_ sg13g2_nand3_1
X_16414_ _08589_ _09235_ _08602_ VPWR VGND _09296_ sg13g2_a21oi_1
X_16415_ _08615_ _09233_ _09294_ _09296_ VPWR VGND 
+ _09297_
+ sg13g2_a22oi_1
X_16416_ _09285_ _09286_ _09295_ _09297_ VPWR VGND 
+ _09298_
+ sg13g2_and4_1
X_16417_ _09165_ _09231_ VPWR VGND _09299_ sg13g2_nand2_1
X_16418_ _09165_ _09231_ _08616_ VPWR VGND _09300_ sg13g2_o21ai_1
X_16419_ _09300_ VPWR VGND _09301_ sg13g2_buf_1
X_16420_ _08456_ _09166_ VPWR VGND _09302_ sg13g2_xor2_1
X_16421_ _08610_ _09302_ VPWR VGND _09303_ sg13g2_nand2_1
X_16422_ _09299_ _09301_ _09303_ VPWR VGND _09304_ sg13g2_a21o_1
X_16423_ _09106_ _09299_ _09301_ _09302_ VPWR VGND 
+ _09305_
+ sg13g2_nand4_1
X_16424_ _08456_ _09166_ VPWR VGND _09306_ sg13g2_xnor2_1
X_16425_ _09106_ _09306_ VPWR VGND _09307_ sg13g2_nand2_1
X_16426_ _09299_ _09301_ _09307_ VPWR VGND _09308_ sg13g2_a21o_1
X_16427_ _08610_ _09299_ _09301_ _09306_ VPWR VGND 
+ _09309_
+ sg13g2_nand4_1
X_16428_ _09304_ _09305_ _09308_ _09309_ VPWR VGND 
+ _09310_
+ sg13g2_nand4_1
X_16429_ _09299_ _09301_ VPWR VGND _09311_ sg13g2_nand2_1
X_16430_ _09311_ _09302_ VPWR VGND _09312_ sg13g2_xnor2_1
X_16431_ _09298_ _09310_ _09312_ _08854_ VPWR VGND 
+ _09313_
+ sg13g2_a22oi_1
X_16432_ _08843_ _09164_ VPWR VGND _09314_ sg13g2_xnor2_1
X_16433_ _09223_ _09314_ VPWR VGND _09315_ sg13g2_xnor2_1
X_16434_ _09229_ _09313_ _09315_ VPWR VGND _09316_ sg13g2_a21oi_1
X_16435_ _09229_ _09313_ VPWR VGND _09317_ sg13g2_nor2_1
X_16436_ _08841_ _09226_ VPWR VGND _09318_ sg13g2_xnor2_1
X_16437_ _09316_ _09317_ _09318_ VPWR VGND _09319_ sg13g2_o21ai_1
X_16438_ _08679_ _09202_ VPWR VGND _09320_ sg13g2_nand2_1
X_16439_ _08940_ _09163_ _09320_ VPWR VGND _09321_ sg13g2_nand3_1
X_16440_ _09202_ _09219_ VPWR VGND _09322_ sg13g2_nand2_1
X_16441_ _09162_ _08704_ VPWR VGND _09323_ sg13g2_xnor2_1
X_16442_ _09321_ _09322_ _09323_ VPWR VGND _09324_ sg13g2_a21oi_1
X_16443_ _08669_ _09163_ _09202_ VPWR VGND _09325_ sg13g2_nor3_1
X_16444_ _08954_ _09203_ _09325_ VPWR VGND _09326_ sg13g2_a21o_1
X_16445_ _09163_ _09202_ _08960_ VPWR VGND _09327_ sg13g2_a21oi_1
X_16446_ _09326_ _09327_ _09323_ VPWR VGND _09328_ sg13g2_o21ai_1
X_16447_ _09324_ _09328_ VPWR VGND _09329_ sg13g2_nor2b_1
X_16448_ _09228_ _09319_ _09329_ VPWR VGND _09330_ sg13g2_a21o_1
X_16449_ _09203_ _09204_ VPWR VGND _09331_ sg13g2_nor2_1
X_16450_ _08726_ _09162_ VPWR VGND _09332_ sg13g2_xor2_1
X_16451_ _09331_ _09332_ VPWR VGND _09333_ sg13g2_xnor2_1
X_16452_ _08729_ _09333_ _08758_ VPWR VGND _09334_ sg13g2_a21oi_1
X_16453_ _09218_ _09330_ _09334_ VPWR VGND _09335_ sg13g2_nand3_1
X_16454_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2656_o[0]\ VPWR VGND _09336_ sg13g2_buf_1
X_16455_ _09336_ VPWR VGND _09337_ sg13g2_inv_1
X_16456_ _09216_ _09335_ _09337_ VPWR VGND _09338_ sg13g2_a21oi_1
X_16457_ _08980_ _09154_ _09338_ VPWR VGND _00498_ sg13g2_a21o_1
X_16458_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2656_o[1]\ VPWR VGND _09339_ sg13g2_buf_1
X_16459_ _09339_ VPWR VGND _09340_ sg13g2_inv_1
X_16460_ _09216_ _09335_ _09340_ VPWR VGND _09341_ sg13g2_a21oi_1
X_16461_ _09150_ _09154_ _09341_ VPWR VGND _00499_ sg13g2_a21o_1
X_16462_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2659_o[0]\ VPWR VGND _09342_ sg13g2_buf_1
X_16463_ _09342_ _09151_ VPWR VGND _09343_ sg13g2_nand2_1
X_16464_ _09336_ _08760_ VPWR VGND _09344_ sg13g2_nand2_1
X_16465_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2661_o\ VPWR VGND _09345_ sg13g2_inv_1
X_16466_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[17]\ VPWR VGND _09346_ sg13g2_buf_1
X_16467_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[16]\ VPWR VGND _09347_ sg13g2_buf_1
X_16468_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[15]\ VPWR VGND _09348_ sg13g2_buf_1
X_16469_ _08667_ _09348_ VPWR VGND _09349_ sg13g2_nor2_1
X_16470_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[13]\ VPWR VGND _09350_ sg13g2_buf_1
X_16471_ _09350_ VPWR VGND _09351_ sg13g2_buf_1
X_16472_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[12]\ VPWR VGND _09352_ sg13g2_buf_1
X_16473_ _08455_ _09352_ VPWR VGND _09353_ sg13g2_nand2_1
X_16474_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[11]\ VPWR VGND _09354_ sg13g2_buf_1
X_16475_ _09354_ VPWR VGND _09355_ sg13g2_inv_1
X_16476_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[9]\ VPWR VGND _09356_ sg13g2_buf_1
X_16477_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[8]\ VPWR VGND _09357_ sg13g2_buf_1
X_16478_ _08416_ _09357_ VPWR VGND _09358_ sg13g2_nor2_1
X_16479_ _09358_ VPWR VGND _09359_ sg13g2_inv_1
X_16480_ _08421_ VPWR VGND _09360_ sg13g2_inv_1
X_16481_ _09360_ VPWR VGND _09361_ sg13g2_buf_2
X_16482_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[6]\ VPWR VGND _09362_ sg13g2_buf_1
X_16483_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[7]\ VPWR VGND _09363_ sg13g2_buf_1
X_16484_ _08424_ _09362_ _09363_ VPWR VGND _09364_ sg13g2_a21oi_1
X_16485_ _08424_ _09363_ _09362_ VPWR VGND _09365_ sg13g2_nand3_1
X_16486_ _09361_ _09364_ _09365_ VPWR VGND _09366_ sg13g2_o21ai_1
X_16487_ _09366_ VPWR VGND _09367_ sg13g2_buf_1
X_16488_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[10]\ VPWR VGND _09368_ sg13g2_buf_1
X_16489_ _08432_ _09368_ _09357_ _08416_ VPWR VGND 
+ _09369_
+ sg13g2_a22oi_1
X_16490_ _09369_ VPWR VGND _09370_ sg13g2_inv_1
X_16491_ _08412_ _09356_ _09359_ _09367_ _09370_ VPWR 
+ VGND
+ _09371_ sg13g2_a221oi_1
X_16492_ _09371_ VPWR VGND _09372_ sg13g2_buf_1
X_16493_ _09356_ VPWR VGND _09373_ sg13g2_inv_1
X_16494_ _08432_ _09368_ VPWR VGND _09374_ sg13g2_nand2_1
X_16495_ _08442_ _09373_ _09374_ VPWR VGND _09375_ sg13g2_nand3_1
X_16496_ _08434_ _09368_ _09375_ VPWR VGND _09376_ sg13g2_o21ai_1
X_16497_ _09355_ _09372_ _09376_ VPWR VGND _09377_ sg13g2_nor3_1
X_16498_ _09372_ _09376_ _09355_ VPWR VGND _09378_ sg13g2_o21ai_1
X_16499_ _08407_ _09377_ _09378_ VPWR VGND _09379_ sg13g2_o21ai_1
X_16500_ _09379_ VPWR VGND _09380_ sg13g2_buf_1
X_16501_ _08456_ _09352_ VPWR VGND _09381_ sg13g2_nor2_1
X_16502_ _09353_ _09380_ _09381_ VPWR VGND _09382_ sg13g2_a21oi_1
X_16503_ _09382_ VPWR VGND _09383_ sg13g2_buf_2
X_16504_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[14]\ VPWR VGND _09384_ sg13g2_buf_1
X_16505_ _09348_ _09384_ VPWR VGND _09385_ sg13g2_or2_1
X_16506_ _08666_ _09384_ VPWR VGND _09386_ sg13g2_or2_1
X_16507_ _09350_ _09352_ _09354_ VPWR VGND _09387_ sg13g2_nor3_1
X_16508_ _08455_ _09350_ _09354_ VPWR VGND _09388_ sg13g2_nor3_1
X_16509_ _09372_ _09376_ VPWR VGND _09389_ sg13g2_or2_1
X_16510_ _09387_ _09388_ _09389_ VPWR VGND _09390_ sg13g2_o21ai_1
X_16511_ _08994_ _09350_ _09352_ VPWR VGND _09391_ sg13g2_nor3_1
X_16512_ _08609_ _08994_ _09351_ VPWR VGND _09392_ sg13g2_nor3_1
X_16513_ _09391_ _09392_ _09389_ VPWR VGND _09393_ sg13g2_o21ai_1
X_16514_ _08609_ _09350_ _09352_ VPWR VGND _09394_ sg13g2_nor3_1
X_16515_ _08407_ _09350_ _09352_ _09354_ VPWR VGND 
+ _09395_
+ sg13g2_nor4_1
X_16516_ _08609_ _08994_ _09350_ _09354_ VPWR VGND 
+ _09396_
+ sg13g2_nor4_1
X_16517_ _09394_ _09395_ _09396_ VPWR VGND _09397_ sg13g2_nor3_1
X_16518_ _08660_ _09390_ _09393_ _09397_ VPWR VGND 
+ _09398_
+ sg13g2_and4_1
X_16519_ _09398_ VPWR VGND _09399_ sg13g2_buf_1
X_16520_ _09351_ _09383_ _09385_ _09386_ _09399_ VPWR 
+ VGND
+ _09400_ sg13g2_a221oi_1
X_16521_ _09348_ VPWR VGND _09401_ sg13g2_inv_1
X_16522_ _08686_ _09401_ VPWR VGND _09402_ sg13g2_nand2_1
X_16523_ _08696_ _08686_ VPWR VGND _09403_ sg13g2_nand2_1
X_16524_ _09351_ _09383_ _09402_ _09403_ _09399_ VPWR 
+ VGND
+ _09404_ sg13g2_a221oi_1
X_16525_ _09402_ _09403_ _09384_ VPWR VGND _09405_ sg13g2_a21oi_1
X_16526_ _09349_ _09400_ _09404_ _09405_ VPWR VGND 
+ _09406_
+ sg13g2_nor4_1
X_16527_ _09347_ _09406_ VPWR VGND _09407_ sg13g2_nand2_1
X_16528_ _09347_ _09406_ _08725_ VPWR VGND _09408_ sg13g2_o21ai_1
X_16529_ _09407_ _09408_ VPWR VGND _09409_ sg13g2_nand2_1
X_16530_ _09346_ _09409_ _08740_ VPWR VGND _09410_ sg13g2_o21ai_1
X_16531_ _09346_ _09409_ VPWR VGND _09411_ sg13g2_nand2_1
X_16532_ _09410_ _09411_ VPWR VGND _09412_ sg13g2_nand2_1
X_16533_ _09384_ VPWR VGND _09413_ sg13g2_buf_1
X_16534_ _09351_ _09383_ _09399_ VPWR VGND _09414_ sg13g2_a21oi_1
X_16535_ _09413_ _09414_ VPWR VGND _09415_ sg13g2_nand2b_1
X_16536_ _09414_ _09413_ VPWR VGND _09416_ sg13g2_nor2b_1
X_16537_ _08682_ _09415_ _09416_ VPWR VGND _09417_ sg13g2_a21oi_1
X_16538_ _08696_ _09401_ VPWR VGND _09418_ sg13g2_nor2_1
X_16539_ _08954_ _09417_ _09418_ VPWR VGND _09419_ sg13g2_o21ai_1
X_16540_ _09347_ _08704_ VPWR VGND _09420_ sg13g2_xnor2_1
X_16541_ _08669_ _09348_ VPWR VGND _09421_ sg13g2_xnor2_1
X_16542_ _09417_ _09421_ VPWR VGND _09422_ sg13g2_nor2_1
X_16543_ _09420_ _09422_ VPWR VGND _09423_ sg13g2_nor2_1
X_16544_ _09413_ _08841_ VPWR VGND _09424_ sg13g2_and2_1
X_16545_ _09413_ _08841_ VPWR VGND _09425_ sg13g2_nor2_1
X_16546_ _09399_ _09424_ _09425_ VPWR VGND _09426_ sg13g2_or3_1
X_16547_ _09351_ _09383_ VPWR VGND _09427_ sg13g2_and2_1
X_16548_ _09394_ _09413_ _08841_ VPWR VGND _09428_ sg13g2_nand3b_1
X_16549_ _09351_ _09383_ _09425_ VPWR VGND _09429_ sg13g2_o21ai_1
X_16550_ _09428_ _09429_ _08849_ VPWR VGND _09430_ sg13g2_a21oi_1
X_16551_ _08849_ _09427_ _09430_ VPWR VGND _09431_ sg13g2_a21oi_1
X_16552_ _09351_ _08676_ _09383_ VPWR VGND _09432_ sg13g2_nand3_1
X_16553_ _09351_ VPWR VGND _09433_ sg13g2_inv_1
X_16554_ _09433_ _08841_ _09353_ _09380_ VPWR VGND 
+ _09434_
+ sg13g2_nand4_1
X_16555_ _09413_ _09432_ _09434_ VPWR VGND _09435_ sg13g2_nand3_1
X_16556_ _08841_ _09427_ _09413_ VPWR VGND _09436_ sg13g2_a21o_1
X_16557_ _09426_ _09431_ _09435_ _09436_ VPWR VGND 
+ _09437_
+ sg13g2_a22oi_1
X_16558_ _08464_ _09351_ VPWR VGND _09438_ sg13g2_xnor2_1
X_16559_ _09383_ _09438_ VPWR VGND _09439_ sg13g2_xnor2_1
X_16560_ _09439_ VPWR VGND _09440_ sg13g2_inv_1
X_16561_ _08570_ _09352_ VPWR VGND _09441_ sg13g2_xnor2_1
X_16562_ _09380_ _09441_ VPWR VGND _09442_ sg13g2_xnor2_1
X_16563_ _08568_ _09442_ VPWR VGND _09443_ sg13g2_nand2_1
X_16564_ _09443_ VPWR VGND _09444_ sg13g2_inv_1
X_16565_ _08551_ _09357_ _09367_ VPWR VGND _09445_ sg13g2_a21oi_1
X_16566_ _09373_ _09358_ _09445_ VPWR VGND _09446_ sg13g2_nor3_1
X_16567_ _09358_ _09445_ _09373_ VPWR VGND _09447_ sg13g2_o21ai_1
X_16568_ _08861_ _09446_ _09447_ VPWR VGND _09448_ sg13g2_o21ai_1
X_16569_ _08595_ _09368_ VPWR VGND _09449_ sg13g2_xnor2_1
X_16570_ _09448_ _09449_ VPWR VGND _09450_ sg13g2_xnor2_1
X_16571_ _09368_ _08623_ VPWR VGND _09451_ sg13g2_xor2_1
X_16572_ _09358_ _09445_ VPWR VGND _09452_ sg13g2_nor2_1
X_16573_ _09356_ _09452_ VPWR VGND _09453_ sg13g2_nor2_1
X_16574_ _08626_ _09446_ _09447_ VPWR VGND _09454_ sg13g2_o21ai_1
X_16575_ _08921_ _09453_ _09454_ _08625_ VPWR VGND 
+ _09455_
+ sg13g2_a22oi_1
X_16576_ _08590_ _09356_ VPWR VGND _09456_ sg13g2_nand2_1
X_16577_ _08626_ _09452_ _09456_ VPWR VGND _09457_ sg13g2_a21oi_1
X_16578_ _08584_ _09356_ VPWR VGND _09458_ sg13g2_xnor2_1
X_16579_ _09358_ _09445_ _09458_ VPWR VGND _09459_ sg13g2_nor3_1
X_16580_ _09457_ _09459_ _09451_ VPWR VGND _09460_ sg13g2_o21ai_1
X_16581_ _09451_ _09455_ _09460_ VPWR VGND _09461_ sg13g2_o21ai_1
X_16582_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ VPWR VGND _09462_ sg13g2_buf_1
X_16583_ _09462_ _08883_ VPWR VGND _09463_ sg13g2_nand2b_1
X_16584_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[154]\ VPWR VGND _09464_ sg13g2_buf_1
X_16585_ _08491_ _09464_ VPWR VGND _09465_ sg13g2_nor2_1
X_16586_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ VPWR VGND _09466_ sg13g2_buf_1
X_16587_ _09466_ _08891_ VPWR VGND _09467_ sg13g2_nand2b_1
X_16588_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ VPWR VGND _09468_ sg13g2_nor2b_1
X_16589_ _08891_ _09466_ VPWR VGND _09469_ sg13g2_nor2b_1
X_16590_ _08491_ _09464_ _09467_ _09468_ _09469_ VPWR 
+ VGND
+ _09470_ sg13g2_a221oi_1
X_16591_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ VPWR VGND _09471_ sg13g2_inv_1
X_16592_ _09465_ _09470_ _09471_ VPWR VGND _09472_ sg13g2_o21ai_1
X_16593_ _09471_ _09465_ _09470_ VPWR VGND _09473_ sg13g2_nor3_1
X_16594_ _08487_ _09472_ _09473_ VPWR VGND _09474_ sg13g2_a21o_1
X_16595_ _08883_ _09462_ VPWR VGND _09475_ sg13g2_nor2b_1
X_16596_ _09463_ _09474_ _09475_ VPWR VGND _09476_ sg13g2_a21oi_1
X_16597_ _08514_ _09362_ VPWR VGND _09477_ sg13g2_nand2_1
X_16598_ _08578_ _09363_ VPWR VGND _09478_ sg13g2_xor2_1
X_16599_ _09477_ _09478_ VPWR VGND _09479_ sg13g2_xnor2_1
X_16600_ _08514_ _09362_ VPWR VGND _09480_ sg13g2_or2_1
X_16601_ _09477_ _09480_ _08907_ VPWR VGND _09481_ sg13g2_a21o_1
X_16602_ _08527_ _09479_ _09481_ VPWR VGND _09482_ sg13g2_o21ai_1
X_16603_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[157]\ VPWR VGND _09483_ sg13g2_buf_1
X_16604_ _09061_ _09483_ VPWR VGND _09484_ sg13g2_nor2_1
X_16605_ _09476_ _09482_ _09484_ VPWR VGND _09485_ sg13g2_nor3_1
X_16606_ _09362_ _08560_ VPWR VGND _09486_ sg13g2_xnor2_1
X_16607_ _09061_ _09483_ _09486_ VPWR VGND _09487_ sg13g2_a21oi_1
X_16608_ _09482_ _09487_ VPWR VGND _09488_ sg13g2_nor2_1
X_16609_ _08872_ _09479_ _09488_ VPWR VGND _09489_ sg13g2_a21oi_1
X_16610_ _08551_ _09357_ VPWR VGND _09490_ sg13g2_xor2_1
X_16611_ _09367_ _09490_ VPWR VGND _09491_ sg13g2_xnor2_1
X_16612_ _08549_ _09491_ VPWR VGND _09492_ sg13g2_xnor2_1
X_16613_ _09489_ _09492_ VPWR VGND _09493_ sg13g2_nand2_1
X_16614_ _09452_ _09458_ VPWR VGND _09494_ sg13g2_xor2_1
X_16615_ _08605_ _09491_ _09494_ _08921_ VPWR VGND 
+ _09495_
+ sg13g2_a22oi_1
X_16616_ _09485_ _09493_ _09495_ VPWR VGND _09496_ sg13g2_o21ai_1
X_16617_ _09048_ _09450_ _09461_ _09496_ VPWR VGND 
+ _09497_
+ sg13g2_a22oi_1
X_16618_ _09377_ _09378_ VPWR VGND _09498_ sg13g2_nand2b_1
X_16619_ _08616_ _09377_ VPWR VGND _09499_ sg13g2_nor2_1
X_16620_ _08617_ _09498_ _09499_ VPWR VGND _09500_ sg13g2_a21oi_1
X_16621_ _08617_ _09378_ VPWR VGND _09501_ sg13g2_nor2_1
X_16622_ _09352_ _08612_ VPWR VGND _09502_ sg13g2_xnor2_1
X_16623_ _09500_ _09501_ _09502_ VPWR VGND _09503_ sg13g2_mux2_1
X_16624_ _08635_ _09503_ VPWR VGND _09504_ sg13g2_nand2_1
X_16625_ _08639_ _09355_ _09502_ VPWR VGND _09505_ sg13g2_nor3_1
X_16626_ _09380_ _09502_ _09505_ VPWR VGND _09506_ sg13g2_a21oi_1
X_16627_ _08615_ _09506_ VPWR VGND _09507_ sg13g2_nor2_1
X_16628_ _09507_ _09503_ VPWR VGND _09508_ sg13g2_nor2_1
X_16629_ _09497_ _09504_ _09508_ VPWR VGND _09509_ sg13g2_a21oi_1
X_16630_ _09440_ _09444_ _09509_ VPWR VGND _09510_ sg13g2_or3_1
X_16631_ _09509_ _09229_ _09443_ VPWR VGND _09511_ sg13g2_nand3b_1
X_16632_ _09229_ _09439_ VPWR VGND _09512_ sg13g2_nand2_1
X_16633_ _09437_ _09510_ _09511_ _09512_ VPWR VGND 
+ _09513_
+ sg13g2_nand4_1
X_16634_ _09417_ _09421_ VPWR VGND _09514_ sg13g2_xnor2_1
X_16635_ _08682_ _09413_ VPWR VGND _09515_ sg13g2_xnor2_1
X_16636_ _09414_ _09515_ VPWR VGND _09516_ sg13g2_xnor2_1
X_16637_ _08954_ _09514_ _09516_ _08943_ VPWR VGND 
+ _09517_
+ sg13g2_a22oi_1
X_16638_ _08679_ _09348_ VPWR VGND _09518_ sg13g2_nor2_1
X_16639_ _09349_ _09518_ _09417_ VPWR VGND _09519_ sg13g2_o21ai_1
X_16640_ _08940_ _08680_ VPWR VGND _09520_ sg13g2_nor2_1
X_16641_ _09401_ _09417_ _09520_ VPWR VGND _09521_ sg13g2_o21ai_1
X_16642_ _09420_ _09519_ _09521_ VPWR VGND _09522_ sg13g2_and3_1
X_16643_ _09419_ _09423_ _09513_ _09517_ _09522_ VPWR 
+ VGND
+ _09523_ sg13g2_a221oi_1
X_16644_ _08726_ _09347_ VPWR VGND _09524_ sg13g2_xnor2_1
X_16645_ _09406_ _09524_ VPWR VGND _09525_ sg13g2_xnor2_1
X_16646_ _09035_ _09525_ VPWR VGND _09526_ sg13g2_nor2_1
X_16647_ _08738_ _09346_ VPWR VGND _09527_ sg13g2_xor2_1
X_16648_ _09409_ _09527_ VPWR VGND _09528_ sg13g2_xnor2_1
X_16649_ _08742_ _09528_ VPWR VGND _09529_ sg13g2_xnor2_1
X_16650_ _09523_ _09526_ _09529_ VPWR VGND _09530_ sg13g2_o21ai_1
X_16651_ _08709_ _09528_ VPWR VGND _09531_ sg13g2_nand2_1
X_16652_ _09345_ _09412_ _09530_ _09531_ _08970_ VPWR 
+ VGND
+ _09532_ sg13g2_a221oi_1
X_16653_ _09343_ _09344_ _09532_ VPWR VGND _00500_ sg13g2_a21oi_1
X_16654_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2659_o[1]\ VPWR VGND _09533_ sg13g2_buf_1
X_16655_ _09533_ VPWR VGND _09534_ sg13g2_buf_1
X_16656_ _09534_ _09151_ VPWR VGND _09535_ sg13g2_nand2_1
X_16657_ _09339_ _08760_ VPWR VGND _09536_ sg13g2_nand2_1
X_16658_ _09535_ _09536_ _09532_ VPWR VGND _00501_ sg13g2_a21oi_1
X_16659_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2662_o[0]\ VPWR VGND _09537_ sg13g2_buf_1
X_16660_ _09537_ _09151_ VPWR VGND _09538_ sg13g2_nand2_1
X_16661_ _09342_ _08760_ VPWR VGND _09539_ sg13g2_nand2_1
X_16662_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[12]\ VPWR VGND _09540_ sg13g2_buf_1
X_16663_ _09540_ _08454_ VPWR VGND _09541_ sg13g2_nand2_1
X_16664_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[14]\ VPWR VGND _09542_ sg13g2_buf_1
X_16665_ _09542_ _08650_ VPWR VGND _09543_ sg13g2_nand2_1
X_16666_ _09541_ _09543_ VPWR VGND _09544_ sg13g2_nand2_1
X_16667_ _08461_ _09544_ VPWR VGND _09545_ sg13g2_nor2_1
X_16668_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[13]\ VPWR VGND _09546_ sg13g2_buf_1
X_16669_ _09546_ _09544_ VPWR VGND _09547_ sg13g2_nor2_1
X_16670_ _09540_ _08609_ VPWR VGND _09548_ sg13g2_or2_1
X_16671_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[9]\ VPWR VGND _09549_ sg13g2_buf_1
X_16672_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[8]\ VPWR VGND _09550_ sg13g2_buf_1
X_16673_ _09550_ _08417_ VPWR VGND _09551_ sg13g2_nor2_1
X_16674_ _09551_ VPWR VGND _09552_ sg13g2_inv_1
X_16675_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[7]\ VPWR VGND _09553_ sg13g2_buf_1
X_16676_ _09553_ VPWR VGND _09554_ sg13g2_inv_1
X_16677_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[6]\ VPWR VGND _09555_ sg13g2_buf_1
X_16678_ _09555_ _08425_ _08422_ VPWR VGND _09556_ sg13g2_a21oi_1
X_16679_ _08422_ _09555_ _08425_ VPWR VGND _09557_ sg13g2_nand3_1
X_16680_ _09554_ _09556_ _09557_ VPWR VGND _09558_ sg13g2_o21ai_1
X_16681_ _09558_ VPWR VGND _09559_ sg13g2_buf_1
X_16682_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[10]\ VPWR VGND _09560_ sg13g2_buf_1
X_16683_ _09560_ _08433_ _09550_ _08417_ VPWR VGND 
+ _09561_
+ sg13g2_a22oi_1
X_16684_ _09561_ VPWR VGND _09562_ sg13g2_inv_1
X_16685_ _09549_ _08412_ _09552_ _09559_ _09562_ VPWR 
+ VGND
+ _09563_ sg13g2_a221oi_1
X_16686_ _09563_ VPWR VGND _09564_ sg13g2_buf_1
X_16687_ _09549_ VPWR VGND _09565_ sg13g2_inv_1
X_16688_ _09560_ _08434_ VPWR VGND _09566_ sg13g2_nand2_1
X_16689_ _09565_ _08443_ _09566_ VPWR VGND _09567_ sg13g2_nand3_1
X_16690_ _09560_ _08441_ _09567_ VPWR VGND _09568_ sg13g2_o21ai_1
X_16691_ _09564_ _09568_ _08638_ VPWR VGND _09569_ sg13g2_o21ai_1
X_16692_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[11]\ VPWR VGND _09570_ sg13g2_inv_1
X_16693_ _09564_ _09568_ _09570_ VPWR VGND _09571_ sg13g2_o21ai_1
X_16694_ _09570_ _08639_ VPWR VGND _09572_ sg13g2_nand2_1
X_16695_ _09548_ _09569_ _09571_ _09572_ VPWR VGND 
+ _09573_
+ sg13g2_nand4_1
X_16696_ _09545_ _09547_ _09573_ VPWR VGND _09574_ sg13g2_o21ai_1
X_16697_ _09546_ _08462_ VPWR VGND _09575_ sg13g2_nor2_1
X_16698_ _09542_ _08651_ VPWR VGND _09576_ sg13g2_nor2_1
X_16699_ _09575_ _09543_ _09576_ VPWR VGND _09577_ sg13g2_a21oi_1
X_16700_ _09574_ _09577_ VPWR VGND _09578_ sg13g2_nand2_1
X_16701_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[15]\ _08669_ VPWR VGND _09579_ sg13g2_xor2_1
X_16702_ _09578_ _09579_ VPWR VGND _09580_ sg13g2_xnor2_1
X_16703_ _09541_ _09573_ VPWR VGND _09581_ sg13g2_nand2_1
X_16704_ _09546_ _08464_ _09581_ VPWR VGND _09582_ sg13g2_a21oi_1
X_16705_ _09575_ _09582_ VPWR VGND _09583_ sg13g2_nor2_1
X_16706_ _09542_ _09583_ VPWR VGND _09584_ sg13g2_xnor2_1
X_16707_ _08841_ _09584_ VPWR VGND _09585_ sg13g2_xnor2_1
X_16708_ _09580_ _09585_ VPWR VGND _09586_ sg13g2_nand2b_1
X_16709_ _08955_ _09585_ VPWR VGND _09587_ sg13g2_nand2_1
X_16710_ _09546_ _08843_ VPWR VGND _09588_ sg13g2_xor2_1
X_16711_ _09581_ _09588_ VPWR VGND _09589_ sg13g2_xnor2_1
X_16712_ _09564_ _09568_ VPWR VGND _09590_ sg13g2_or2_1
X_16713_ _08639_ _09590_ _09570_ VPWR VGND _09591_ sg13g2_o21ai_1
X_16714_ _09591_ _09569_ VPWR VGND _09592_ sg13g2_nand2_1
X_16715_ _09540_ _08570_ VPWR VGND _09593_ sg13g2_xnor2_1
X_16716_ _09592_ _09593_ VPWR VGND _09594_ sg13g2_xnor2_1
X_16717_ _08854_ _09594_ VPWR VGND _09595_ sg13g2_nand2_1
X_16718_ _09550_ _08550_ VPWR VGND _09596_ sg13g2_and2_1
X_16719_ _09552_ _09559_ _09596_ VPWR VGND _09597_ sg13g2_a21o_1
X_16720_ _09597_ VPWR VGND _09598_ sg13g2_buf_1
X_16721_ _09549_ _08583_ VPWR VGND _09599_ sg13g2_xor2_1
X_16722_ _09549_ _08590_ VPWR VGND _09600_ sg13g2_nand2_1
X_16723_ _08626_ _09598_ _09600_ VPWR VGND _09601_ sg13g2_a21oi_1
X_16724_ _09598_ _09599_ _09601_ VPWR VGND _09602_ sg13g2_a21oi_1
X_16725_ _09560_ _08623_ VPWR VGND _09603_ sg13g2_xor2_1
X_16726_ _08576_ _09598_ VPWR VGND _09604_ sg13g2_nor2_1
X_16727_ _08626_ _09598_ _08590_ VPWR VGND _09605_ sg13g2_a21oi_1
X_16728_ _09604_ _09605_ _09565_ VPWR VGND _09606_ sg13g2_o21ai_1
X_16729_ _08625_ _09604_ _09603_ VPWR VGND _09607_ sg13g2_a21oi_1
X_16730_ _09602_ _09603_ _09606_ _09607_ VPWR VGND 
+ _09608_
+ sg13g2_a22oi_1
X_16731_ _09553_ _08868_ VPWR VGND _09609_ sg13g2_xor2_1
X_16732_ _09555_ _08514_ VPWR VGND _09610_ sg13g2_and2_1
X_16733_ _09610_ VPWR VGND _09611_ sg13g2_buf_1
X_16734_ _09550_ _08436_ VPWR VGND _09612_ sg13g2_xnor2_1
X_16735_ _08548_ _09612_ VPWR VGND _09613_ sg13g2_xor2_1
X_16736_ _09613_ VPWR VGND _09614_ sg13g2_buf_1
X_16737_ _09614_ _08534_ VPWR VGND _09615_ sg13g2_nand2b_1
X_16738_ _08872_ _09611_ _09614_ VPWR VGND _09616_ sg13g2_nand3_1
X_16739_ _09611_ _09615_ _09616_ VPWR VGND _09617_ sg13g2_o21ai_1
X_16740_ _08534_ _09611_ VPWR VGND _09618_ sg13g2_xnor2_1
X_16741_ _08868_ _09614_ _09554_ VPWR VGND _09619_ sg13g2_a21oi_1
X_16742_ _08868_ _09614_ _09554_ VPWR VGND _09620_ sg13g2_o21ai_1
X_16743_ _09619_ _09620_ VPWR VGND _09621_ sg13g2_nor2b_1
X_16744_ _09609_ _09617_ _09618_ _09621_ VPWR VGND 
+ _09622_
+ sg13g2_a22oi_1
X_16745_ _09555_ _08542_ VPWR VGND _09623_ sg13g2_xor2_1
X_16746_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[176]\ VPWR VGND _09624_ sg13g2_buf_1
X_16747_ _08508_ _09624_ _09061_ VPWR VGND _09625_ sg13g2_nor3_1
X_16748_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ VPWR VGND _09626_ sg13g2_buf_1
X_16749_ _09626_ _08882_ VPWR VGND _09627_ sg13g2_nand2b_1
X_16750_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ VPWR VGND _09628_ sg13g2_buf_1
X_16751_ _09628_ _08889_ VPWR VGND _09629_ sg13g2_nor2_1
X_16752_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[172]\ VPWR VGND _09630_ sg13g2_buf_1
X_16753_ _09630_ _08891_ VPWR VGND _09631_ sg13g2_nand2b_1
X_16754_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ VPWR VGND _09632_ sg13g2_nor2b_1
X_16755_ _09071_ _09630_ VPWR VGND _09633_ sg13g2_nor2b_1
X_16756_ _09628_ _08491_ _09631_ _09632_ _09633_ VPWR 
+ VGND
+ _09634_ sg13g2_a221oi_1
X_16757_ _09629_ _09634_ _08885_ VPWR VGND _09635_ sg13g2_o21ai_1
X_16758_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _09627_ _09635_ VPWR VGND _09636_ sg13g2_nand3_1
X_16759_ _09555_ _08560_ VPWR VGND _09637_ sg13g2_xnor2_1
X_16760_ _08882_ _09626_ VPWR VGND _09638_ sg13g2_nor2b_1
X_16761_ _09624_ _08878_ VPWR VGND _09639_ sg13g2_xor2_1
X_16762_ _08487_ _09627_ VPWR VGND _09640_ sg13g2_nand2_1
X_16763_ _09629_ _09634_ _09640_ VPWR VGND _09641_ sg13g2_nor3_1
X_16764_ _09637_ _09638_ _09639_ _09641_ VPWR VGND 
+ _09642_
+ sg13g2_nor4_1
X_16765_ _09624_ _08878_ _08508_ VPWR VGND _09643_ sg13g2_nand3b_1
X_16766_ _08907_ _09643_ _09623_ VPWR VGND _09644_ sg13g2_a21oi_1
X_16767_ _09623_ _09625_ _09636_ _09642_ _09644_ VPWR 
+ VGND
+ _09645_ sg13g2_a221oi_1
X_16768_ _09559_ _09612_ VPWR VGND _09646_ sg13g2_xor2_1
X_16769_ _09598_ _09599_ VPWR VGND _09647_ sg13g2_xnor2_1
X_16770_ _09554_ _09557_ VPWR VGND _09648_ sg13g2_nand2_1
X_16771_ _08867_ _09555_ _08514_ VPWR VGND _09649_ sg13g2_and3_1
X_16772_ _09556_ _09649_ _09553_ VPWR VGND _09650_ sg13g2_o21ai_1
X_16773_ _09648_ _09614_ _09650_ VPWR VGND _09651_ sg13g2_nand3_1
X_16774_ _09553_ _08868_ _09611_ _09614_ VPWR VGND 
+ _09652_
+ sg13g2_or4_1
X_16775_ _09651_ _09652_ _08872_ VPWR VGND _09653_ sg13g2_a21oi_1
X_16776_ _08604_ _09646_ _09647_ _08920_ _09653_ VPWR 
+ VGND
+ _09654_ sg13g2_a221oi_1
X_16777_ _09622_ _09645_ _09654_ VPWR VGND _09655_ sg13g2_o21ai_1
X_16778_ _08590_ _09598_ _09549_ VPWR VGND _09656_ sg13g2_a21oi_1
X_16779_ _08590_ _09598_ VPWR VGND _09657_ sg13g2_nor2_1
X_16780_ _09656_ _09657_ VPWR VGND _09658_ sg13g2_nor2_1
X_16781_ _09560_ _08595_ VPWR VGND _09659_ sg13g2_xor2_1
X_16782_ _09658_ _09659_ VPWR VGND _09660_ sg13g2_xnor2_1
X_16783_ _09608_ _09655_ _09660_ _09048_ VPWR VGND 
+ _09661_
+ sg13g2_a22oi_1
X_16784_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[11]\ _08617_ VPWR VGND _09662_ sg13g2_xor2_1
X_16785_ _09590_ _09662_ VPWR VGND _09663_ sg13g2_xnor2_1
X_16786_ _08930_ _09661_ _09663_ VPWR VGND _09664_ sg13g2_a21oi_1
X_16787_ _08930_ _09661_ VPWR VGND _09665_ sg13g2_nor2_1
X_16788_ _08610_ _09594_ VPWR VGND _09666_ sg13g2_xnor2_1
X_16789_ _09664_ _09665_ _09666_ VPWR VGND _09667_ sg13g2_o21ai_1
X_16790_ _09229_ _09595_ _09667_ VPWR VGND _09668_ sg13g2_nand3_1
X_16791_ _09595_ _09667_ _09229_ VPWR VGND _09669_ sg13g2_a21oi_1
X_16792_ _09589_ _09668_ _09669_ VPWR VGND _09670_ sg13g2_a21oi_1
X_16793_ _09586_ _09587_ _09670_ VPWR VGND _09671_ sg13g2_a21oi_1
X_16794_ _08685_ _08687_ _09584_ VPWR VGND _09672_ sg13g2_mux2_1
X_16795_ _08681_ _09580_ _09672_ VPWR VGND _09673_ sg13g2_a21o_1
X_16796_ _08681_ _09580_ _09673_ VPWR VGND _09674_ sg13g2_o21ai_1
X_16797_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[16]\ VPWR VGND _09675_ sg13g2_buf_1
X_16798_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[15]\ VPWR VGND _09676_ sg13g2_inv_1
X_16799_ _08666_ _09574_ _09577_ VPWR VGND _09677_ sg13g2_nand3_1
X_16800_ _09574_ _09577_ _08667_ VPWR VGND _09678_ sg13g2_a21oi_1
X_16801_ _09676_ _09677_ _09678_ VPWR VGND _09679_ sg13g2_a21oi_1
X_16802_ _09675_ _09679_ VPWR VGND _09680_ sg13g2_xor2_1
X_16803_ _08704_ _09680_ VPWR VGND _09681_ sg13g2_xnor2_1
X_16804_ _09671_ _09674_ _09681_ VPWR VGND _09682_ sg13g2_o21ai_1
X_16805_ _08726_ _09680_ VPWR VGND _09683_ sg13g2_xnor2_1
X_16806_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[17]\ VPWR VGND _09684_ sg13g2_buf_1
X_16807_ _09675_ _08701_ VPWR VGND _09685_ sg13g2_and2_1
X_16808_ _09675_ _08701_ VPWR VGND _09686_ sg13g2_or2_1
X_16809_ _09685_ _09679_ _09686_ VPWR VGND _09687_ sg13g2_o21ai_1
X_16810_ _09687_ VPWR VGND _09688_ sg13g2_buf_1
X_16811_ _08738_ _09688_ VPWR VGND _09689_ sg13g2_xnor2_1
X_16812_ _09684_ _09689_ VPWR VGND _09690_ sg13g2_xnor2_1
X_16813_ _08729_ _09683_ _09690_ _08709_ VPWR VGND 
+ _09691_
+ sg13g2_a22oi_1
X_16814_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2664_o\ VPWR VGND _09692_ sg13g2_buf_1
X_16815_ _08711_ _09688_ VPWR VGND _09693_ sg13g2_nor2_1
X_16816_ _09693_ _09689_ _09684_ VPWR VGND _09694_ sg13g2_mux2_1
X_16817_ _08712_ _09688_ VPWR VGND _09695_ sg13g2_nand2_1
X_16818_ _09684_ _09695_ _08741_ VPWR VGND _09696_ sg13g2_o21ai_1
X_16819_ _09692_ _09694_ _09696_ VPWR VGND _09697_ sg13g2_a21o_1
X_16820_ _08708_ _09689_ VPWR VGND _09698_ sg13g2_nor2_1
X_16821_ _08712_ _09692_ _09688_ VPWR VGND _09699_ sg13g2_nor3_1
X_16822_ _09684_ _08741_ VPWR VGND _09700_ sg13g2_nor2_1
X_16823_ _09698_ _09699_ _09700_ VPWR VGND _09701_ sg13g2_o21ai_1
X_16824_ _08708_ _09693_ _09692_ VPWR VGND _09702_ sg13g2_o21ai_1
X_16825_ _09684_ _08744_ _09695_ _09702_ VPWR VGND 
+ _09703_
+ sg13g2_nand4_1
X_16826_ _07931_ _09697_ _09701_ _09703_ VPWR VGND 
+ _09704_
+ sg13g2_nand4_1
X_16827_ _09682_ _09691_ _09704_ VPWR VGND _09705_ sg13g2_a21oi_1
X_16828_ _09538_ _09539_ _09705_ VPWR VGND _00502_ sg13g2_a21oi_1
X_16829_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2662_o[1]\ VPWR VGND _09706_ sg13g2_buf_1
X_16830_ _09706_ _09151_ VPWR VGND _09707_ sg13g2_nand2_1
X_16831_ _09534_ _08760_ VPWR VGND _09708_ sg13g2_nand2_1
X_16832_ _09707_ _09708_ _09705_ VPWR VGND _00503_ sg13g2_a21oi_1
X_16833_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2635_o[1]\ VPWR VGND _09709_ sg13g2_buf_1
X_16834_ _09709_ VPWR VGND _09710_ sg13g2_inv_1
X_16835_ _08754_ _07799_ VPWR VGND _09711_ sg13g2_nor2b_1
X_16836_ _09710_ _07799_ _08731_ _09711_ _07733_ VPWR 
+ VGND
+ _00504_ sg13g2_a221oi_1
X_16837_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2665_o[0]\ VPWR VGND _09712_ sg13g2_buf_1
X_16838_ _09712_ _09151_ VPWR VGND _09713_ sg13g2_nand2_1
X_16839_ _09537_ _08760_ VPWR VGND _09714_ sg13g2_nand2_1
X_16840_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[15]\ VPWR VGND _09715_ sg13g2_buf_1
X_16841_ _08667_ _09715_ VPWR VGND _09716_ sg13g2_xor2_1
X_16842_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[14]\ VPWR VGND _09717_ sg13g2_buf_1
X_16843_ _08675_ _09717_ VPWR VGND _09718_ sg13g2_nand2_1
X_16844_ _09716_ _09718_ VPWR VGND _09719_ sg13g2_nor2_1
X_16845_ _08675_ VPWR VGND _09720_ sg13g2_buf_1
X_16846_ _08667_ _09715_ VPWR VGND _09721_ sg13g2_xnor2_1
X_16847_ _09720_ _09717_ _09721_ VPWR VGND _09722_ sg13g2_nor3_1
X_16848_ _09719_ _09722_ _08679_ VPWR VGND _09723_ sg13g2_o21ai_1
X_16849_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[11]\ VPWR VGND _09724_ sg13g2_buf_1
X_16850_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[10]\ VPWR VGND _09725_ sg13g2_buf_1
X_16851_ _08594_ _09725_ VPWR VGND _09726_ sg13g2_or2_1
X_16852_ _09726_ VPWR VGND _09727_ sg13g2_buf_1
X_16853_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[8]\ VPWR VGND _09728_ sg13g2_buf_1
X_16854_ _08417_ _09728_ VPWR VGND _09729_ sg13g2_nor2_1
X_16855_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[6]\ VPWR VGND _09730_ sg13g2_buf_2
X_16856_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[7]\ VPWR VGND _09731_ sg13g2_buf_1
X_16857_ _08423_ _09730_ _09731_ VPWR VGND _09732_ sg13g2_a21o_1
X_16858_ _09732_ VPWR VGND _09733_ sg13g2_buf_1
X_16859_ _08424_ _09731_ _09730_ VPWR VGND _09734_ sg13g2_and3_1
X_16860_ _09734_ VPWR VGND _09735_ sg13g2_buf_1
X_16861_ _08416_ _09728_ _09733_ _08422_ _09735_ VPWR 
+ VGND
+ _09736_ sg13g2_a221oi_1
X_16862_ _09736_ VPWR VGND _09737_ sg13g2_buf_1
X_16863_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[9]\ VPWR VGND _09738_ sg13g2_buf_1
X_16864_ _09738_ VPWR VGND _09739_ sg13g2_inv_1
X_16865_ _09729_ _09737_ _09739_ VPWR VGND _09740_ sg13g2_o21ai_1
X_16866_ _09740_ VPWR VGND _09741_ sg13g2_buf_1
X_16867_ _09739_ _09729_ _09737_ VPWR VGND _09742_ sg13g2_nor3_1
X_16868_ _08413_ _09741_ _09742_ VPWR VGND _09743_ sg13g2_a21o_1
X_16869_ _09743_ VPWR VGND _09744_ sg13g2_buf_1
X_16870_ _08594_ _09725_ VPWR VGND _09745_ sg13g2_and2_1
X_16871_ _09745_ VPWR VGND _09746_ sg13g2_buf_1
X_16872_ _08994_ _09724_ _09727_ _09744_ _09746_ VPWR 
+ VGND
+ _09747_ sg13g2_a221oi_1
X_16873_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[12]\ VPWR VGND _09748_ sg13g2_buf_1
X_16874_ _08453_ _09748_ VPWR VGND _09749_ sg13g2_or2_1
X_16875_ _09749_ VPWR VGND _09750_ sg13g2_buf_1
X_16876_ _08408_ _09724_ _09750_ VPWR VGND _09751_ sg13g2_o21ai_1
X_16877_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[13]\ VPWR VGND _09752_ sg13g2_buf_1
X_16878_ _08456_ _09748_ _09752_ VPWR VGND _09753_ sg13g2_a21oi_1
X_16879_ _09747_ _09751_ _09753_ VPWR VGND _09754_ sg13g2_o21ai_1
X_16880_ _08594_ _09725_ VPWR VGND _09755_ sg13g2_nor2_1
X_16881_ _08594_ _09725_ _09741_ _08413_ _09742_ VPWR 
+ VGND
+ _09756_ sg13g2_a221oi_1
X_16882_ _09756_ VPWR VGND _09757_ sg13g2_buf_1
X_16883_ _09752_ _09724_ _09750_ VPWR VGND _09758_ sg13g2_nand3_1
X_16884_ _09755_ _09757_ _09758_ VPWR VGND _09759_ sg13g2_nor3_1
X_16885_ _08407_ _09752_ _09750_ VPWR VGND _09760_ sg13g2_nand3_1
X_16886_ _09755_ _09757_ _09760_ VPWR VGND _09761_ sg13g2_nor3_1
X_16887_ _09724_ VPWR VGND _09762_ sg13g2_inv_1
X_16888_ _08455_ _09752_ _09748_ VPWR VGND _09763_ sg13g2_nand3_1
X_16889_ _09762_ _09760_ _09763_ VPWR VGND _09764_ sg13g2_o21ai_1
X_16890_ _08462_ _09759_ _09761_ _09764_ VPWR VGND 
+ _09765_
+ sg13g2_or4_1
X_16891_ _09754_ _09765_ VPWR VGND _09766_ sg13g2_and2_1
X_16892_ _09766_ VPWR VGND _09767_ sg13g2_buf_1
X_16893_ _08675_ _09717_ VPWR VGND _09768_ sg13g2_xnor2_1
X_16894_ _09767_ _09768_ VPWR VGND _09769_ sg13g2_xnor2_1
X_16895_ _08679_ _09716_ _09718_ VPWR VGND _09770_ sg13g2_nand3_1
X_16896_ _09769_ _09770_ _08682_ VPWR VGND _09771_ sg13g2_a21o_1
X_16897_ _08675_ _09717_ _08679_ VPWR VGND _09772_ sg13g2_o21ai_1
X_16898_ _09716_ _09772_ VPWR VGND _09773_ sg13g2_nor2_1
X_16899_ _09769_ _09773_ _08682_ VPWR VGND _09774_ sg13g2_o21ai_1
X_16900_ _09755_ _09746_ VPWR VGND _09775_ sg13g2_nor2_1
X_16901_ _09744_ _09775_ VPWR VGND _09776_ sg13g2_xnor2_1
X_16902_ _09725_ _08622_ VPWR VGND _09777_ sg13g2_xor2_1
X_16903_ _08575_ _09742_ _09741_ VPWR VGND _09778_ sg13g2_o21ai_1
X_16904_ _08575_ _09741_ VPWR VGND _09779_ sg13g2_nor2_1
X_16905_ _08443_ _09778_ _09779_ VPWR VGND _09780_ sg13g2_a21oi_1
X_16906_ _08413_ _09738_ VPWR VGND _09781_ sg13g2_xnor2_1
X_16907_ _09729_ _09737_ _09781_ VPWR VGND _09782_ sg13g2_nor3_1
X_16908_ _09729_ _09737_ VPWR VGND _09783_ sg13g2_nor2_1
X_16909_ _08583_ _09738_ VPWR VGND _09784_ sg13g2_nand2_1
X_16910_ _08575_ _09783_ _09784_ VPWR VGND _09785_ sg13g2_a21oi_1
X_16911_ _09782_ _09785_ _09777_ VPWR VGND _09786_ sg13g2_o21ai_1
X_16912_ _09777_ _09780_ _09786_ VPWR VGND _09787_ sg13g2_o21ai_1
X_16913_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ VPWR VGND _09788_ sg13g2_inv_1
X_16914_ _09730_ _08560_ VPWR VGND _09789_ sg13g2_xnor2_1
X_16915_ _09733_ VPWR VGND _09790_ sg13g2_inv_1
X_16916_ _08468_ _09735_ _09733_ VPWR VGND _09791_ sg13g2_o21ai_1
X_16917_ _08416_ _08548_ VPWR VGND _09792_ sg13g2_xor2_1
X_16918_ _09728_ _09792_ VPWR VGND _09793_ sg13g2_xnor2_1
X_16919_ _08532_ _09790_ _09791_ _09361_ _09793_ VPWR 
+ VGND
+ _09794_ sg13g2_a221oi_1
X_16920_ _08469_ _09731_ VPWR VGND _09795_ sg13g2_and2_1
X_16921_ _08513_ _08468_ _09730_ VPWR VGND _09796_ sg13g2_nand3_1
X_16922_ _08469_ _09731_ VPWR VGND _09797_ sg13g2_xor2_1
X_16923_ _08513_ _09730_ VPWR VGND _09798_ sg13g2_and2_1
X_16924_ _09795_ _09796_ _09797_ _09798_ VPWR VGND 
+ _09799_
+ sg13g2_a22oi_1
X_16925_ _09793_ _09799_ VPWR VGND _09800_ sg13g2_and2_1
X_16926_ _09789_ _09794_ _09800_ VPWR VGND _09801_ sg13g2_nor3_1
X_16927_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[193]\ VPWR VGND _09802_ sg13g2_inv_1
X_16928_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ VPWR VGND _09803_ sg13g2_inv_1
X_16929_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[191]\ VPWR VGND _09804_ sg13g2_buf_1
X_16930_ _09804_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[1]\ VPWR VGND _09805_ sg13g2_nand2b_1
X_16931_ _08494_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ VPWR VGND _09806_ sg13g2_nor2b_1
X_16932_ _08498_ _09804_ VPWR VGND _09807_ sg13g2_nor2b_1
X_16933_ _08490_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ _09805_ _09806_ _09807_ VPWR 
+ VGND
+ _09808_ sg13g2_a221oi_1
X_16934_ _08485_ _09802_ _09803_ _08489_ _09808_ VPWR 
+ VGND
+ _09809_ sg13g2_a221oi_1
X_16935_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ VPWR VGND _09810_ sg13g2_buf_1
X_16936_ _08482_ _09810_ VPWR VGND _09811_ sg13g2_nand2_1
X_16937_ _08485_ _09802_ _09811_ VPWR VGND _09812_ sg13g2_o21ai_1
X_16938_ _09810_ _08882_ VPWR VGND _09813_ sg13g2_nand2b_1
X_16939_ _09809_ _09812_ _09813_ VPWR VGND _09814_ sg13g2_o21ai_1
X_16940_ _09788_ _09801_ _09814_ VPWR VGND _09815_ sg13g2_nand3_1
X_16941_ _08477_ _09789_ _09794_ _09800_ VPWR VGND 
+ _09816_
+ sg13g2_nor4_1
X_16942_ _09788_ _09814_ _09816_ VPWR VGND _09817_ sg13g2_o21ai_1
X_16943_ _09783_ _09781_ VPWR VGND _09818_ sg13g2_nor2b_1
X_16944_ _09782_ _09818_ _08920_ VPWR VGND _09819_ sg13g2_o21ai_1
X_16945_ _08513_ _09731_ _09730_ VPWR VGND _09820_ sg13g2_nand3_1
X_16946_ _09733_ _09820_ _09361_ VPWR VGND _09821_ sg13g2_a21oi_1
X_16947_ _09361_ _09820_ _09821_ VPWR VGND _09822_ sg13g2_a21oi_1
X_16948_ _08867_ _09733_ _09793_ VPWR VGND _09823_ sg13g2_nor3_1
X_16949_ _09793_ _09822_ _09823_ VPWR VGND _09824_ sg13g2_a21o_1
X_16950_ _08513_ _09730_ VPWR VGND _09825_ sg13g2_nor2_1
X_16951_ _09798_ _09825_ _08555_ VPWR VGND _09826_ sg13g2_o21ai_1
X_16952_ _08527_ _09826_ VPWR VGND _09827_ sg13g2_nand2_1
X_16953_ _08527_ _09826_ VPWR VGND _09828_ sg13g2_nor2_1
X_16954_ _08578_ _09733_ _09735_ VPWR VGND _09829_ sg13g2_a21oi_1
X_16955_ _09829_ _09795_ _09793_ VPWR VGND _09830_ sg13g2_mux2_1
X_16956_ _08550_ _09728_ VPWR VGND _09831_ sg13g2_xnor2_1
X_16957_ _09829_ _09831_ VPWR VGND _09832_ sg13g2_xnor2_1
X_16958_ _08604_ _09832_ VPWR VGND _09833_ sg13g2_and2_1
X_16959_ _09824_ _09827_ _09828_ _09830_ _09833_ VPWR 
+ VGND
+ _09834_ sg13g2_a221oi_1
X_16960_ _09815_ _09817_ _09819_ _09834_ VPWR VGND 
+ _09835_
+ sg13g2_nand4_1
X_16961_ _09755_ _09757_ VPWR VGND _09836_ sg13g2_nor2_1
X_16962_ _08408_ _09724_ VPWR VGND _09837_ sg13g2_xor2_1
X_16963_ _09836_ _09837_ VPWR VGND _09838_ sg13g2_xnor2_1
X_16964_ _08589_ _09776_ _09787_ _09835_ _09838_ VPWR 
+ VGND
+ _09839_ sg13g2_a221oi_1
X_16965_ _08589_ _09776_ _09787_ _09835_ _08635_ VPWR 
+ VGND
+ _09840_ sg13g2_a221oi_1
X_16966_ _08635_ _09838_ VPWR VGND _09841_ sg13g2_nor2_1
X_16967_ _09839_ _09840_ _09841_ VPWR VGND _09842_ sg13g2_nor3_1
X_16968_ _09757_ _09724_ _09727_ VPWR VGND _09843_ sg13g2_nand3b_1
X_16969_ _09724_ _09746_ VPWR VGND _09844_ sg13g2_nor2_1
X_16970_ _09727_ _09744_ VPWR VGND _09845_ sg13g2_nand2_1
X_16971_ _08639_ _09843_ _09844_ _09845_ VPWR VGND 
+ _09846_
+ sg13g2_a22oi_1
X_16972_ _09846_ VPWR VGND _09847_ sg13g2_buf_1
X_16973_ _08455_ _09748_ VPWR VGND _09848_ sg13g2_xnor2_1
X_16974_ _09106_ _09847_ _09848_ VPWR VGND _09849_ sg13g2_nor3_1
X_16975_ _08610_ _09848_ VPWR VGND _09850_ sg13g2_nor2_1
X_16976_ _09847_ _09850_ VPWR VGND _09851_ sg13g2_and2_1
X_16977_ _09106_ _09848_ VPWR VGND _09852_ sg13g2_and2_1
X_16978_ _08610_ _09848_ VPWR VGND _09853_ sg13g2_and2_1
X_16979_ _09852_ _09853_ _09847_ VPWR VGND _09854_ sg13g2_mux2_1
X_16980_ _09849_ _09851_ _09854_ VPWR VGND _09855_ sg13g2_nor3_1
X_16981_ _09847_ _09848_ VPWR VGND _09856_ sg13g2_xnor2_1
X_16982_ _08570_ _09748_ VPWR VGND _09857_ sg13g2_nand2_1
X_16983_ _09747_ _09751_ _09857_ VPWR VGND _09858_ sg13g2_o21ai_1
X_16984_ _08463_ _09752_ VPWR VGND _09859_ sg13g2_xnor2_1
X_16985_ _09858_ _09859_ VPWR VGND _09860_ sg13g2_xnor2_1
X_16986_ _08569_ _09856_ _09860_ VPWR VGND _09861_ sg13g2_o21ai_1
X_16987_ _09842_ _09855_ _09861_ VPWR VGND _09862_ sg13g2_a21o_1
X_16988_ _09723_ _09771_ _09774_ _09862_ VPWR VGND 
+ _09863_
+ sg13g2_and4_1
X_16989_ _08569_ _09856_ VPWR VGND _09864_ sg13g2_nor2_1
X_16990_ _09842_ _09855_ _09864_ VPWR VGND _09865_ sg13g2_a21oi_1
X_16991_ _09860_ _09865_ _09229_ VPWR VGND _09866_ sg13g2_o21ai_1
X_16992_ _08682_ _09717_ VPWR VGND _09867_ sg13g2_xnor2_1
X_16993_ _08683_ VPWR VGND _09868_ sg13g2_inv_1
X_16994_ _09767_ _09867_ _09868_ VPWR VGND _09869_ sg13g2_a21oi_1
X_16995_ _09869_ _08680_ VPWR VGND _09870_ sg13g2_nand2b_1
X_16996_ _09868_ _09767_ _08679_ VPWR VGND _09871_ sg13g2_a21oi_1
X_16997_ _08653_ _09717_ VPWR VGND _09872_ sg13g2_or2_1
X_16998_ _09872_ VPWR VGND _09873_ sg13g2_buf_1
X_16999_ _09721_ _09873_ VPWR VGND _09874_ sg13g2_nand2_1
X_17000_ _09871_ _09874_ VPWR VGND _09875_ sg13g2_nor2_1
X_17001_ _08679_ _09868_ _09767_ VPWR VGND _09876_ sg13g2_nor3_1
X_17002_ _09721_ _09873_ _09876_ VPWR VGND _09877_ sg13g2_nor3_1
X_17003_ _09868_ _09767_ VPWR VGND _09878_ sg13g2_or2_1
X_17004_ _08653_ _09717_ VPWR VGND _09879_ sg13g2_and2_1
X_17005_ _09721_ _09878_ _09879_ VPWR VGND _09880_ sg13g2_and3_1
X_17006_ _09721_ _09767_ _09867_ VPWR VGND _09881_ sg13g2_nor3_1
X_17007_ _09875_ _09877_ _09880_ _09881_ VPWR VGND 
+ _09882_
+ sg13g2_nor4_1
X_17008_ _09863_ _09866_ _09870_ _09882_ VPWR VGND 
+ _09883_
+ sg13g2_a22oi_1
X_17009_ _08668_ _09715_ VPWR VGND _09884_ sg13g2_nand2_1
X_17010_ _09767_ _09879_ _09873_ VPWR VGND _09885_ sg13g2_o21ai_1
X_17011_ _08668_ _09715_ VPWR VGND _09886_ sg13g2_nor2_1
X_17012_ _09884_ _09885_ _09886_ VPWR VGND _09887_ sg13g2_a21oi_1
X_17013_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[16]\ VPWR VGND _09888_ sg13g2_buf_1
X_17014_ _09205_ _09888_ VPWR VGND _09889_ sg13g2_xnor2_1
X_17015_ _09887_ _09889_ VPWR VGND _09890_ sg13g2_xnor2_1
X_17016_ _08702_ _09890_ VPWR VGND _09891_ sg13g2_xnor2_1
X_17017_ _09035_ _09890_ VPWR VGND _09892_ sg13g2_or2_1
X_17018_ _09883_ _09891_ _09892_ VPWR VGND _09893_ sg13g2_o21ai_1
X_17019_ _08742_ _09893_ _08709_ VPWR VGND _09894_ sg13g2_a21oi_1
X_17020_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2667_o\ VPWR VGND _09895_ sg13g2_inv_1
X_17021_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[17]\ VPWR VGND _09896_ sg13g2_buf_1
X_17022_ _09205_ _09888_ VPWR VGND _09897_ sg13g2_and2_1
X_17023_ _09897_ VPWR VGND _09898_ sg13g2_buf_1
X_17024_ _09896_ _09898_ _08739_ VPWR VGND _09899_ sg13g2_o21ai_1
X_17025_ _09896_ _09898_ VPWR VGND _09900_ sg13g2_nand2_1
X_17026_ _09899_ _09900_ VPWR VGND _09901_ sg13g2_nand2_1
X_17027_ _08725_ _09888_ VPWR VGND _09902_ sg13g2_or2_1
X_17028_ _08739_ _09896_ _09902_ VPWR VGND _09903_ sg13g2_o21ai_1
X_17029_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2667_o\ _09903_ VPWR VGND _09904_ sg13g2_nor2_1
X_17030_ _09895_ _09901_ _09904_ _09887_ _08758_ VPWR 
+ VGND
+ _09905_ sg13g2_a221oi_1
X_17031_ _08739_ _09896_ VPWR VGND _09906_ sg13g2_xnor2_1
X_17032_ _09887_ _09902_ _09898_ VPWR VGND _09907_ sg13g2_a21oi_1
X_17033_ _09906_ _09907_ VPWR VGND _09908_ sg13g2_xnor2_1
X_17034_ _09905_ _09908_ VPWR VGND _09909_ sg13g2_nand2_1
X_17035_ _08742_ _09908_ VPWR VGND _09910_ sg13g2_nor2_1
X_17036_ _09893_ _09905_ _09910_ VPWR VGND _09911_ sg13g2_nand3_1
X_17037_ _09894_ _09909_ _09911_ VPWR VGND _09912_ sg13g2_o21ai_1
X_17038_ _09713_ _09714_ _09912_ VPWR VGND _00505_ sg13g2_a21oi_1
X_17039_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2665_o[1]\ VPWR VGND _09913_ sg13g2_buf_1
X_17040_ _09913_ VPWR VGND _09914_ sg13g2_buf_1
X_17041_ _09914_ _09151_ VPWR VGND _09915_ sg13g2_nand2_1
X_17042_ _09706_ _08981_ VPWR VGND _09916_ sg13g2_nand2_1
X_17043_ _09915_ _09916_ _09912_ VPWR VGND _00506_ sg13g2_a21oi_1
X_17044_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[12]\ VPWR VGND _09917_ sg13g2_buf_1
X_17045_ _09917_ VPWR VGND _09918_ sg13g2_inv_1
X_17046_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[11]\ VPWR VGND _09919_ sg13g2_buf_1
X_17047_ _08994_ _09919_ VPWR VGND _09920_ sg13g2_nor2_1
X_17048_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[8]\ VPWR VGND _09921_ sg13g2_buf_1
X_17049_ _08416_ _09921_ VPWR VGND _09922_ sg13g2_nor2_1
X_17050_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[6]\ VPWR VGND _09923_ sg13g2_buf_1
X_17051_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[7]\ VPWR VGND _09924_ sg13g2_buf_1
X_17052_ _08424_ _09923_ _09924_ VPWR VGND _09925_ sg13g2_a21o_1
X_17053_ _08424_ _09924_ _09923_ VPWR VGND _09926_ sg13g2_and3_1
X_17054_ _08415_ _09921_ _09925_ _08421_ _09926_ VPWR 
+ VGND
+ _09927_ sg13g2_a221oi_1
X_17055_ _09927_ VPWR VGND _09928_ sg13g2_buf_1
X_17056_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[9]\ VPWR VGND _09929_ sg13g2_buf_1
X_17057_ _09929_ VPWR VGND _09930_ sg13g2_inv_1
X_17058_ _09922_ _09928_ _09930_ VPWR VGND _09931_ sg13g2_o21ai_1
X_17059_ _09931_ VPWR VGND _09932_ sg13g2_buf_1
X_17060_ _09930_ _09922_ _09928_ VPWR VGND _09933_ sg13g2_nor3_1
X_17061_ _08413_ _09932_ _09933_ VPWR VGND _09934_ sg13g2_a21o_1
X_17062_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[10]\ VPWR VGND _09935_ sg13g2_buf_1
X_17063_ _08441_ _09935_ VPWR VGND _09936_ sg13g2_nor2_1
X_17064_ _09936_ VPWR VGND _09937_ sg13g2_inv_1
X_17065_ _08441_ VPWR VGND _09938_ sg13g2_inv_1
X_17066_ _09935_ VPWR VGND _09939_ sg13g2_inv_1
X_17067_ _09938_ _09939_ VPWR VGND _09940_ sg13g2_nor2_1
X_17068_ _08407_ _09919_ _09934_ _09937_ _09940_ VPWR 
+ VGND
+ _09941_ sg13g2_a221oi_1
X_17069_ _09918_ _09920_ _09941_ VPWR VGND _09942_ sg13g2_nor3_1
X_17070_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[13]\ VPWR VGND _09943_ sg13g2_buf_1
X_17071_ _08461_ _09943_ VPWR VGND _09944_ sg13g2_or2_1
X_17072_ _09944_ VPWR VGND _09945_ sg13g2_buf_1
X_17073_ _09942_ _09945_ VPWR VGND _09946_ sg13g2_nand2_1
X_17074_ _08441_ _09935_ VPWR VGND _09947_ sg13g2_nand2_1
X_17075_ _09917_ _09919_ VPWR VGND _09948_ sg13g2_nor2_1
X_17076_ _09947_ _09948_ VPWR VGND _09949_ sg13g2_nand2_1
X_17077_ _08405_ _09917_ VPWR VGND _09950_ sg13g2_nor2_1
X_17078_ _09947_ _09950_ VPWR VGND _09951_ sg13g2_nand2_1
X_17079_ _08413_ _09932_ _09949_ _09951_ _09933_ VPWR 
+ VGND
+ _09952_ sg13g2_a221oi_1
X_17080_ _09952_ VPWR VGND _09953_ sg13g2_buf_1
X_17081_ _08406_ _09917_ _09919_ VPWR VGND _09954_ sg13g2_nor3_1
X_17082_ _09948_ _09950_ _09936_ VPWR VGND _09955_ sg13g2_o21ai_1
X_17083_ _09954_ _09955_ VPWR VGND _09956_ sg13g2_nand2b_1
X_17084_ _09956_ VPWR VGND _09957_ sg13g2_buf_1
X_17085_ _09953_ _09957_ VPWR VGND _09958_ sg13g2_nor2_1
X_17086_ _08570_ _09958_ _09945_ VPWR VGND _09959_ sg13g2_nand3_1
X_17087_ _08461_ _09943_ VPWR VGND _09960_ sg13g2_nand2_1
X_17088_ _09960_ VPWR VGND _09961_ sg13g2_buf_1
X_17089_ _08686_ _09946_ _09959_ _09961_ VPWR VGND 
+ _09962_
+ sg13g2_nand4_1
X_17090_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[14]\ VPWR VGND _09963_ sg13g2_buf_1
X_17091_ _09963_ VPWR VGND _09964_ sg13g2_inv_1
X_17092_ _09964_ _09946_ _09959_ _09961_ VPWR VGND 
+ _09965_
+ sg13g2_nand4_1
X_17093_ _08686_ _09964_ VPWR VGND _09966_ sg13g2_nand2_1
X_17094_ _09962_ _09965_ _09966_ VPWR VGND _09967_ sg13g2_nand3_1
X_17095_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[15]\ VPWR VGND _09968_ sg13g2_buf_1
X_17096_ _08669_ _09968_ VPWR VGND _09969_ sg13g2_xnor2_1
X_17097_ _09967_ _09969_ VPWR VGND _09970_ sg13g2_xnor2_1
X_17098_ _09963_ _08676_ VPWR VGND _09971_ sg13g2_xnor2_1
X_17099_ _09961_ _09971_ VPWR VGND _09972_ sg13g2_nor2_1
X_17100_ _08462_ _09943_ VPWR VGND _09973_ sg13g2_xnor2_1
X_17101_ _09971_ _09973_ VPWR VGND _09974_ sg13g2_nor2_1
X_17102_ _08787_ _09971_ _09973_ VPWR VGND _09975_ sg13g2_nor3_1
X_17103_ _09942_ _09974_ _09975_ _09958_ VPWR VGND 
+ _09976_
+ sg13g2_a22oi_1
X_17104_ _09917_ _09919_ VPWR VGND _09977_ sg13g2_nand2_1
X_17105_ _08406_ _09917_ VPWR VGND _09978_ sg13g2_nand2_1
X_17106_ _08582_ _09932_ _09933_ VPWR VGND _09979_ sg13g2_a21oi_1
X_17107_ _09938_ _09939_ _09977_ _09978_ _09979_ VPWR 
+ VGND
+ _09980_ sg13g2_a221oi_1
X_17108_ _09980_ VPWR VGND _09981_ sg13g2_buf_1
X_17109_ _09977_ _09978_ _09947_ VPWR VGND _09982_ sg13g2_a21oi_1
X_17110_ _08408_ _09917_ _09919_ VPWR VGND _09983_ sg13g2_nand3_1
X_17111_ _09982_ _09983_ VPWR VGND _09984_ sg13g2_nand2b_1
X_17112_ _09981_ _09984_ VPWR VGND _09985_ sg13g2_nor2_1
X_17113_ _08461_ _09943_ VPWR VGND _09986_ sg13g2_nor2_1
X_17114_ _09986_ _09971_ _09972_ VPWR VGND _09987_ sg13g2_a21o_1
X_17115_ _08787_ _09987_ VPWR VGND _09988_ sg13g2_and2_1
X_17116_ _09958_ _09987_ VPWR VGND _09989_ sg13g2_nor2b_1
X_17117_ _09985_ _09988_ _09989_ VPWR VGND _09990_ sg13g2_a21oi_1
X_17118_ _09976_ _09990_ VPWR VGND _09991_ sg13g2_nand2_1
X_17119_ _09946_ _09959_ _09961_ _09971_ VPWR VGND 
+ _09992_
+ sg13g2_and4_1
X_17120_ _08650_ _09963_ VPWR VGND _09993_ sg13g2_xnor2_1
X_17121_ _09993_ _08683_ _09945_ VPWR VGND _09994_ sg13g2_nand3b_1
X_17122_ _08787_ _09953_ _09957_ _09994_ VPWR VGND 
+ _09995_
+ sg13g2_nor4_1
X_17123_ _08787_ _09953_ _09957_ VPWR VGND _09996_ sg13g2_nor3_1
X_17124_ _08683_ _09961_ _09993_ VPWR VGND _09997_ sg13g2_nand3_1
X_17125_ _09981_ _09984_ _09996_ _09997_ VPWR VGND 
+ _09998_
+ sg13g2_nor4_1
X_17126_ _09918_ _09920_ _09941_ _09994_ VPWR VGND 
+ _09999_
+ sg13g2_nor4_1
X_17127_ _08660_ _08683_ _09943_ VPWR VGND _10000_ sg13g2_nand3_1
X_17128_ _08683_ _09986_ _09993_ VPWR VGND _10001_ sg13g2_nand3_1
X_17129_ _09993_ _10000_ _10001_ VPWR VGND _10002_ sg13g2_o21ai_1
X_17130_ _09995_ _09998_ _09999_ _10002_ VPWR VGND 
+ _10003_
+ sg13g2_or4_1
X_17131_ _09972_ _09991_ _09992_ _10003_ VPWR VGND 
+ _10004_
+ sg13g2_nor4_1
X_17132_ _09979_ _09936_ _09947_ VPWR VGND _10005_ sg13g2_o21ai_1
X_17133_ _08616_ _09919_ VPWR VGND _10006_ sg13g2_xnor2_1
X_17134_ _10005_ _10006_ VPWR VGND _10007_ sg13g2_xnor2_1
X_17135_ _09940_ _09936_ VPWR VGND _10008_ sg13g2_nor2_1
X_17136_ _09934_ _10008_ VPWR VGND _10009_ sg13g2_xnor2_1
X_17137_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ VPWR VGND _10010_ sg13g2_inv_1
X_17138_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ VPWR VGND _10011_ sg13g2_inv_1
X_17139_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ VPWR VGND _10012_ sg13g2_buf_1
X_17140_ _10012_ _08489_ VPWR VGND _10013_ sg13g2_nand2b_1
X_17141_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ VPWR VGND _10014_ sg13g2_buf_1
X_17142_ _10014_ _08498_ VPWR VGND _10015_ sg13g2_nor2b_1
X_17143_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ VPWR VGND _10016_ sg13g2_nand2b_1
X_17144_ _08891_ _10014_ VPWR VGND _10017_ sg13g2_nand2b_1
X_17145_ _10015_ _10016_ _10017_ VPWR VGND _10018_ sg13g2_o21ai_1
X_17146_ _08888_ _10012_ VPWR VGND _10019_ sg13g2_nor2b_1
X_17147_ _08486_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _10013_ _10018_ _10019_ VPWR 
+ VGND
+ _10020_ sg13g2_a221oi_1
X_17148_ _08885_ _10010_ _10011_ _08882_ _10020_ VPWR 
+ VGND
+ _10021_ sg13g2_a221oi_1
X_17149_ _08883_ _10011_ VPWR VGND _10022_ sg13g2_nor2_1
X_17150_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ VPWR VGND _10023_ sg13g2_inv_1
X_17151_ _08514_ _09923_ VPWR VGND _10024_ sg13g2_xnor2_1
X_17152_ _08878_ _10023_ _10024_ _08556_ VPWR VGND 
+ _10025_
+ sg13g2_a22oi_1
X_17153_ _10021_ _10022_ _10025_ VPWR VGND _10026_ sg13g2_o21ai_1
X_17154_ _08477_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ VPWR VGND _10027_ sg13g2_nand2_1
X_17155_ _08508_ _10027_ _08556_ VPWR VGND _10028_ sg13g2_a21oi_1
X_17156_ _08542_ _09923_ VPWR VGND _10029_ sg13g2_nand2_1
X_17157_ _08867_ _09924_ VPWR VGND _10030_ sg13g2_xor2_1
X_17158_ _10029_ _10030_ VPWR VGND _10031_ sg13g2_xnor2_1
X_17159_ _08475_ _10027_ _10024_ VPWR VGND _10032_ sg13g2_a21oi_1
X_17160_ _10024_ _10028_ _10031_ _08872_ _10032_ VPWR 
+ VGND
+ _10033_ sg13g2_a221oi_1
X_17161_ _08872_ _10031_ VPWR VGND _10034_ sg13g2_nor2_1
X_17162_ _10026_ _10033_ _10034_ VPWR VGND _10035_ sg13g2_a21o_1
X_17163_ _09935_ _08622_ VPWR VGND _10036_ sg13g2_xnor2_1
X_17164_ _09922_ _09928_ VPWR VGND _10037_ sg13g2_nor2_1
X_17165_ _08583_ _09929_ VPWR VGND _10038_ sg13g2_nand2_1
X_17166_ _08575_ _10037_ _10038_ VPWR VGND _10039_ sg13g2_a21oi_1
X_17167_ _08582_ _09929_ VPWR VGND _10040_ sg13g2_xnor2_1
X_17168_ _09922_ _09928_ _10040_ VPWR VGND _10041_ sg13g2_nor3_1
X_17169_ _10036_ _10039_ _10041_ VPWR VGND _10042_ sg13g2_nor3_1
X_17170_ _08575_ _09932_ VPWR VGND _10043_ sg13g2_nor2_1
X_17171_ _08413_ _08574_ VPWR VGND _10044_ sg13g2_nor2_1
X_17172_ _09933_ _10044_ VPWR VGND _10045_ sg13g2_nor2b_1
X_17173_ _08584_ _09932_ _10036_ VPWR VGND _10046_ sg13g2_o21ai_1
X_17174_ _10043_ _10045_ _10046_ VPWR VGND _10047_ sg13g2_nor3_1
X_17175_ _08867_ _09925_ _09926_ VPWR VGND _10048_ sg13g2_a21oi_1
X_17176_ _08550_ _09921_ VPWR VGND _10049_ sg13g2_xnor2_1
X_17177_ _10048_ _10049_ VPWR VGND _10050_ sg13g2_xnor2_1
X_17178_ _08549_ _10050_ VPWR VGND _10051_ sg13g2_xor2_1
X_17179_ _10042_ _10047_ _10051_ VPWR VGND _10052_ sg13g2_nor3_1
X_17180_ _10037_ _10040_ VPWR VGND _10053_ sg13g2_xor2_1
X_17181_ _08604_ _10050_ _10053_ _08920_ VPWR VGND 
+ _10054_
+ sg13g2_a22oi_1
X_17182_ _10042_ _10047_ _10054_ VPWR VGND _10055_ sg13g2_nor3_1
X_17183_ _08589_ _10009_ _10035_ _10052_ _10055_ VPWR 
+ VGND
+ _10056_ sg13g2_a221oi_1
X_17184_ _08615_ _10007_ _10056_ VPWR VGND _10057_ sg13g2_o21ai_1
X_17185_ _09981_ _09984_ _09953_ _09957_ VPWR VGND 
+ _10058_
+ sg13g2_nor4_1
X_17186_ _08612_ _10058_ VPWR VGND _10059_ sg13g2_nand2b_1
X_17187_ _10058_ _08612_ VPWR VGND _10060_ sg13g2_nand2b_1
X_17188_ _08615_ _10007_ VPWR VGND _10061_ sg13g2_nand2_1
X_17189_ _10059_ _10060_ _10061_ VPWR VGND _10062_ sg13g2_and3_1
X_17190_ _08787_ _08568_ VPWR VGND _10063_ sg13g2_nand2_1
X_17191_ _08570_ _08568_ VPWR VGND _10064_ sg13g2_nand2_1
X_17192_ _10063_ _10064_ _10058_ VPWR VGND _10065_ sg13g2_mux2_1
X_17193_ _09995_ _09998_ _09999_ _10002_ VPWR VGND 
+ _10066_
+ sg13g2_nor4_1
X_17194_ _09976_ _09990_ _10065_ _10066_ VPWR VGND 
+ _10067_
+ sg13g2_nand4_1
X_17195_ _10057_ _10062_ _10067_ VPWR VGND _10068_ sg13g2_a21oi_1
X_17196_ _08644_ _10065_ _10066_ VPWR VGND _10069_ sg13g2_nand3_1
X_17197_ _10057_ _10062_ _10069_ VPWR VGND _10070_ sg13g2_a21oi_1
X_17198_ _08646_ _09991_ _10003_ VPWR VGND _10071_ sg13g2_nor3_1
X_17199_ _10004_ _10068_ _10070_ _10071_ VPWR VGND 
+ _10072_
+ sg13g2_nor4_1
X_17200_ _09970_ _10072_ _08955_ VPWR VGND _10073_ sg13g2_o21ai_1
X_17201_ _09970_ _10072_ VPWR VGND _10074_ sg13g2_nand2_1
X_17202_ _10073_ _10074_ VPWR VGND _10075_ sg13g2_nand2_1
X_17203_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[16]\ VPWR VGND _10076_ sg13g2_buf_1
X_17204_ _08666_ _09968_ VPWR VGND _10077_ sg13g2_nor2_1
X_17205_ _08666_ _09968_ VPWR VGND _10078_ sg13g2_nand2_1
X_17206_ _09964_ _09961_ _10078_ VPWR VGND _10079_ sg13g2_nand3_1
X_17207_ _08686_ _09961_ _10078_ VPWR VGND _10080_ sg13g2_nand3_1
X_17208_ _08787_ _09953_ _09957_ _09986_ VPWR VGND 
+ _10081_
+ sg13g2_nor4_1
X_17209_ _09942_ _09945_ _10079_ _10080_ _10081_ VPWR 
+ VGND
+ _10082_ sg13g2_a221oi_1
X_17210_ _09966_ _10078_ VPWR VGND _10083_ sg13g2_nor2b_1
X_17211_ _10077_ _10082_ _10083_ VPWR VGND _10084_ sg13g2_nor3_1
X_17212_ _10076_ _10084_ VPWR VGND _10085_ sg13g2_xnor2_1
X_17213_ _08704_ _10085_ VPWR VGND _10086_ sg13g2_xor2_1
X_17214_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[17]\ VPWR VGND _10087_ sg13g2_buf_1
X_17215_ _08724_ _10076_ _10084_ VPWR VGND _10088_ sg13g2_a21o_1
X_17216_ _09205_ _10076_ _10088_ VPWR VGND _10089_ sg13g2_o21ai_1
X_17217_ _10089_ VPWR VGND _10090_ sg13g2_buf_1
X_17218_ _10087_ _10090_ VPWR VGND _10091_ sg13g2_xnor2_1
X_17219_ _08822_ _10091_ VPWR VGND _10092_ sg13g2_xnor2_1
X_17220_ _08726_ _10085_ VPWR VGND _10093_ sg13g2_xnor2_1
X_17221_ _09035_ _10093_ VPWR VGND _10094_ sg13g2_nor2_1
X_17222_ _10075_ _10086_ _10092_ _08708_ _10094_ VPWR 
+ VGND
+ _10095_ sg13g2_a221oi_1
X_17223_ _08822_ _10087_ VPWR VGND _10096_ sg13g2_nor2_1
X_17224_ _10087_ VPWR VGND _10097_ sg13g2_inv_1
X_17225_ _08739_ _10097_ _10090_ VPWR VGND _10098_ sg13g2_nor3_1
X_17226_ _08822_ _10091_ _10098_ VPWR VGND _10099_ sg13g2_a21o_1
X_17227_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2670_o\ VPWR VGND _10100_ sg13g2_buf_1
X_17228_ _10090_ _10096_ _10099_ _10100_ _08744_ VPWR 
+ VGND
+ _10101_ sg13g2_a221oi_1
X_17229_ _08822_ _10087_ _10100_ VPWR VGND _10102_ sg13g2_nand3_1
X_17230_ _08822_ _10097_ _10090_ VPWR VGND _10103_ sg13g2_nand3_1
X_17231_ _10090_ _10102_ _10103_ VPWR VGND _10104_ sg13g2_o21ai_1
X_17232_ _08707_ _10087_ VPWR VGND _10105_ sg13g2_nor2_1
X_17233_ _10087_ _10105_ _10090_ VPWR VGND _10106_ sg13g2_mux2_1
X_17234_ _08708_ _10100_ _08741_ VPWR VGND _10107_ sg13g2_a21oi_1
X_17235_ _08740_ _10106_ _10107_ VPWR VGND _10108_ sg13g2_o21ai_1
X_17236_ _10104_ _10108_ _07931_ VPWR VGND _10109_ sg13g2_o21ai_1
X_17237_ _10095_ _10101_ _10109_ VPWR VGND _10110_ sg13g2_nor3_1
X_17238_ _09712_ _09151_ VPWR VGND _10111_ sg13g2_nor2_1
X_17239_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2668_o[0]\ VPWR VGND _10112_ sg13g2_buf_1
X_17240_ _10112_ _08760_ VPWR VGND _10113_ sg13g2_nor2_1
X_17241_ _10110_ _10111_ _10113_ VPWR VGND _00507_ sg13g2_nor3_1
X_17242_ _09914_ _08977_ VPWR VGND _10114_ sg13g2_nor2_1
X_17243_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2668_o[1]\ VPWR VGND _10115_ sg13g2_buf_1
X_17244_ _10115_ _08760_ VPWR VGND _10116_ sg13g2_nor2_1
X_17245_ _10110_ _10114_ _10116_ VPWR VGND _00508_ sg13g2_nor3_1
X_17246_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[16]\ VPWR VGND _10117_ sg13g2_buf_1
X_17247_ _08724_ _10117_ VPWR VGND _10118_ sg13g2_nor2_1
X_17248_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[12]\ VPWR VGND _10119_ sg13g2_buf_1
X_17249_ _08609_ _10119_ VPWR VGND _10120_ sg13g2_nor2_1
X_17250_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[10]\ VPWR VGND _10121_ sg13g2_buf_1
X_17251_ _08432_ _10121_ VPWR VGND _10122_ sg13g2_nand2_1
X_17252_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[9]\ VPWR VGND _10123_ sg13g2_buf_1
X_17253_ _08415_ VPWR VGND _10124_ sg13g2_inv_1
X_17254_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[8]\ VPWR VGND _10125_ sg13g2_buf_1
X_17255_ _10125_ VPWR VGND _10126_ sg13g2_inv_1
X_17256_ _10124_ _10126_ VPWR VGND _10127_ sg13g2_nor2_1
X_17257_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[7]\ VPWR VGND _10128_ sg13g2_buf_1
X_17258_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[6]\ VPWR VGND _10129_ sg13g2_buf_2
X_17259_ _08424_ _10128_ _10129_ VPWR VGND _10130_ sg13g2_nand3_1
X_17260_ _08424_ _10129_ _10128_ VPWR VGND _10131_ sg13g2_a21oi_1
X_17261_ _09361_ _10130_ _10131_ VPWR VGND _10132_ sg13g2_a21oi_1
X_17262_ _10123_ VPWR VGND _10133_ sg13g2_inv_1
X_17263_ _10124_ _10126_ _10133_ VPWR VGND _10134_ sg13g2_a21oi_1
X_17264_ _10123_ _10127_ _10132_ _10134_ _08412_ VPWR 
+ VGND
+ _10135_ sg13g2_a221oi_1
X_17265_ _10124_ _10126_ _10130_ _09361_ _10131_ VPWR 
+ VGND
+ _10136_ sg13g2_a221oi_1
X_17266_ _10136_ VPWR VGND _10137_ sg13g2_buf_1
X_17267_ _08416_ _10125_ VPWR VGND _10138_ sg13g2_nand2_1
X_17268_ _10133_ _10122_ _10138_ VPWR VGND _10139_ sg13g2_nand3_1
X_17269_ _08433_ _10121_ VPWR VGND _10140_ sg13g2_or2_1
X_17270_ _10137_ _10139_ _10140_ VPWR VGND _10141_ sg13g2_o21ai_1
X_17271_ _10122_ _10135_ _10141_ VPWR VGND _10142_ sg13g2_a21oi_1
X_17272_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[11]\ VPWR VGND _10143_ sg13g2_buf_1
X_17273_ _08405_ _10143_ VPWR VGND _10144_ sg13g2_or2_1
X_17274_ _08405_ _10143_ VPWR VGND _10145_ sg13g2_and2_1
X_17275_ _08454_ _10119_ _10142_ _10144_ _10145_ VPWR 
+ VGND
+ _10146_ sg13g2_a221oi_1
X_17276_ _10146_ VPWR VGND _10147_ sg13g2_buf_1
X_17277_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[13]\ VPWR VGND _10148_ sg13g2_inv_1
X_17278_ _10120_ _10147_ _10148_ VPWR VGND _10149_ sg13g2_o21ai_1
X_17279_ _08455_ _10119_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[13]\ VPWR VGND _10150_ sg13g2_o21ai_1
X_17280_ _10147_ _10150_ _08848_ VPWR VGND _10151_ sg13g2_o21ai_1
X_17281_ _10149_ _10151_ VPWR VGND _10152_ sg13g2_nand2_1
X_17282_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[14]\ VPWR VGND _10153_ sg13g2_buf_1
X_17283_ _08652_ _10153_ VPWR VGND _10154_ sg13g2_nand2_1
X_17284_ _08652_ _10153_ VPWR VGND _10155_ sg13g2_nor2_1
X_17285_ _10152_ _10154_ _10155_ VPWR VGND _10156_ sg13g2_a21oi_1
X_17286_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[15]\ VPWR VGND _10157_ sg13g2_buf_1
X_17287_ _08667_ _10157_ VPWR VGND _10158_ sg13g2_and2_1
X_17288_ _08667_ _10157_ VPWR VGND _10159_ sg13g2_or2_1
X_17289_ _10156_ _10158_ _10159_ VPWR VGND _10160_ sg13g2_o21ai_1
X_17290_ _09205_ _10117_ VPWR VGND _10161_ sg13g2_nand2_1
X_17291_ _10118_ _10160_ _10161_ VPWR VGND _10162_ sg13g2_o21ai_1
X_17292_ _10162_ VPWR VGND _10163_ sg13g2_buf_1
X_17293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[17]\ VPWR VGND _10164_ sg13g2_buf_1
X_17294_ _08738_ _10164_ VPWR VGND _10165_ sg13g2_xor2_1
X_17295_ _10163_ _10165_ VPWR VGND _10166_ sg13g2_xnor2_1
X_17296_ _10166_ _08744_ VPWR VGND _10167_ sg13g2_nand2b_1
X_17297_ _08742_ _10166_ VPWR VGND _10168_ sg13g2_nand2_1
X_17298_ _08725_ _10117_ VPWR VGND _10169_ sg13g2_xnor2_1
X_17299_ _10160_ _10169_ VPWR VGND _10170_ sg13g2_xnor2_1
X_17300_ _08702_ _10170_ VPWR VGND _10171_ sg13g2_xnor2_1
X_17301_ _08668_ _10157_ VPWR VGND _10172_ sg13g2_xor2_1
X_17302_ _10156_ _10172_ VPWR VGND _10173_ sg13g2_xnor2_1
X_17303_ _10155_ _10154_ VPWR VGND _10174_ sg13g2_nor2b_1
X_17304_ _10152_ _10174_ VPWR VGND _10175_ sg13g2_xnor2_1
X_17305_ _09868_ _10175_ VPWR VGND _10176_ sg13g2_nor2_1
X_17306_ _08954_ _10173_ _10176_ VPWR VGND _10177_ sg13g2_o21ai_1
X_17307_ _10142_ _10144_ _10145_ VPWR VGND _10178_ sg13g2_a21oi_1
X_17308_ _08456_ _10119_ VPWR VGND _10179_ sg13g2_xnor2_1
X_17309_ _10178_ _10179_ VPWR VGND _10180_ sg13g2_xnor2_1
X_17310_ _08610_ _10180_ VPWR VGND _10181_ sg13g2_xnor2_1
X_17311_ _10127_ _10137_ VPWR VGND _10182_ sg13g2_nor2_1
X_17312_ _10133_ _10182_ _10135_ VPWR VGND _10183_ sg13g2_a21oi_1
X_17313_ _10122_ _10140_ VPWR VGND _10184_ sg13g2_and2_1
X_17314_ _10183_ _10184_ VPWR VGND _10185_ sg13g2_xnor2_1
X_17315_ _08550_ _10125_ VPWR VGND _10186_ sg13g2_xor2_1
X_17316_ _10132_ _10186_ VPWR VGND _10187_ sg13g2_xnor2_1
X_17317_ _08549_ _10187_ VPWR VGND _10188_ sg13g2_xor2_1
X_17318_ _08469_ _10128_ VPWR VGND _10189_ sg13g2_xor2_1
X_17319_ _08527_ _10189_ VPWR VGND _10190_ sg13g2_nand2_1
X_17320_ _10129_ _10190_ VPWR VGND _10191_ sg13g2_nor2_1
X_17321_ _09270_ VPWR VGND _10192_ sg13g2_buf_1
X_17322_ _08533_ _10192_ VPWR VGND _10193_ sg13g2_nor2_1
X_17323_ _08533_ _10192_ _10189_ VPWR VGND _10194_ sg13g2_a21oi_1
X_17324_ _10193_ _10194_ _10129_ VPWR VGND _10195_ sg13g2_o21ai_1
X_17325_ _10129_ VPWR VGND _10196_ sg13g2_inv_1
X_17326_ _10189_ _08532_ VPWR VGND _10197_ sg13g2_nand2b_1
X_17327_ _10197_ VPWR VGND _10198_ sg13g2_buf_1
X_17328_ _08508_ _10196_ _10198_ VPWR VGND _10199_ sg13g2_nand3_1
X_17329_ _10195_ _10199_ _08516_ VPWR VGND _10200_ sg13g2_a21oi_1
X_17330_ _08474_ _10129_ VPWR VGND _10201_ sg13g2_nand2_1
X_17331_ _10129_ _10192_ _10201_ VPWR VGND _10202_ sg13g2_o21ai_1
X_17332_ _10198_ _10202_ VPWR VGND _10203_ sg13g2_nand2_1
X_17333_ _10190_ _10203_ _08543_ VPWR VGND _10204_ sg13g2_a21oi_1
X_17334_ _10188_ _10191_ _10200_ _10204_ VPWR VGND 
+ _10205_
+ sg13g2_nor4_1
X_17335_ _10121_ _08622_ VPWR VGND _10206_ sg13g2_xor2_1
X_17336_ _10127_ _10137_ VPWR VGND _10207_ sg13g2_or2_1
X_17337_ _08582_ _10123_ VPWR VGND _10208_ sg13g2_xor2_1
X_17338_ _08443_ _10133_ VPWR VGND _10209_ sg13g2_nor2_1
X_17339_ _10127_ _10137_ _08575_ VPWR VGND _10210_ sg13g2_o21ai_1
X_17340_ _10207_ _10208_ _10209_ _10210_ VPWR VGND 
+ _10211_
+ sg13g2_a22oi_1
X_17341_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[233]\ VPWR VGND _10212_ sg13g2_buf_1
X_17342_ _08476_ _10212_ VPWR VGND _10213_ sg13g2_nor2b_1
X_17343_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ VPWR VGND _10214_ sg13g2_buf_1
X_17344_ _08882_ _10214_ VPWR VGND _10215_ sg13g2_nor2b_1
X_17345_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ VPWR VGND _10216_ sg13g2_inv_1
X_17346_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[229]\ VPWR VGND _10217_ sg13g2_buf_1
X_17347_ _09071_ _10217_ VPWR VGND _10218_ sg13g2_nand2b_1
X_17348_ _10217_ _08891_ VPWR VGND _10219_ sg13g2_nand2b_1
X_17349_ _08894_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ _10219_ VPWR VGND _10220_ sg13g2_nand3b_1
X_17350_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ VPWR VGND _10221_ sg13g2_buf_1
X_17351_ _08889_ _10221_ VPWR VGND _10222_ sg13g2_nor2_1
X_17352_ _08485_ _10216_ _10218_ _10220_ _10222_ VPWR 
+ VGND
+ _10223_ sg13g2_a221oi_1
X_17353_ _08489_ _10221_ VPWR VGND _10224_ sg13g2_nor2b_1
X_17354_ _08486_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ _10224_ VPWR VGND _10225_ sg13g2_o21ai_1
X_17355_ _08485_ _10216_ _10225_ VPWR VGND _10226_ sg13g2_o21ai_1
X_17356_ _10213_ _10215_ _10223_ _10226_ VPWR VGND 
+ _10227_
+ sg13g2_or4_1
X_17357_ _08533_ _10189_ _08556_ VPWR VGND _10228_ sg13g2_a21oi_1
X_17358_ _08515_ _10196_ _10228_ VPWR VGND _10229_ sg13g2_nor3_1
X_17359_ _08556_ _10196_ VPWR VGND _10230_ sg13g2_nand2_1
X_17360_ _10198_ _10230_ _08542_ VPWR VGND _10231_ sg13g2_a21oi_1
X_17361_ _10129_ _10198_ VPWR VGND _10232_ sg13g2_nor2_1
X_17362_ _10214_ _08480_ VPWR VGND _10233_ sg13g2_nand2b_1
X_17363_ _10212_ _10233_ _08477_ VPWR VGND _10234_ sg13g2_o21ai_1
X_17364_ _10212_ _10233_ VPWR VGND _10235_ sg13g2_nand2_1
X_17365_ _10234_ _10235_ VPWR VGND _10236_ sg13g2_and2_1
X_17366_ _10229_ _10231_ _10232_ _10236_ VPWR VGND 
+ _10237_
+ sg13g2_nor4_1
X_17367_ _08443_ _10133_ VPWR VGND _10238_ sg13g2_nand2_1
X_17368_ _08920_ _10133_ VPWR VGND _10239_ sg13g2_nand2_1
X_17369_ _08551_ _10125_ _10238_ _10239_ _10137_ VPWR 
+ VGND
+ _10240_ sg13g2_a221oi_1
X_17370_ _08583_ _08575_ _10127_ _10137_ VPWR VGND 
+ _10241_
+ sg13g2_nor4_1
X_17371_ _08583_ _08575_ _10123_ VPWR VGND _10242_ sg13g2_nor3_1
X_17372_ _10206_ _10240_ _10241_ _10242_ VPWR VGND 
+ _10243_
+ sg13g2_nor4_1
X_17373_ _10206_ _10211_ _10227_ _10237_ _10243_ VPWR 
+ VGND
+ _10244_ sg13g2_a221oi_1
X_17374_ _08920_ _10208_ VPWR VGND _10245_ sg13g2_and2_1
X_17375_ _08604_ _10187_ _10245_ _10207_ VPWR VGND 
+ _10246_
+ sg13g2_a22oi_1
X_17376_ _10208_ _08920_ _10182_ VPWR VGND _10247_ sg13g2_nand3b_1
X_17377_ _10206_ _10211_ _10246_ _10247_ _10243_ VPWR 
+ VGND
+ _10248_ sg13g2_a221oi_1
X_17378_ _08589_ _10185_ _10205_ _10244_ _10248_ VPWR 
+ VGND
+ _10249_ sg13g2_a221oi_1
X_17379_ _08617_ _10143_ VPWR VGND _10250_ sg13g2_xnor2_1
X_17380_ _10142_ _10250_ VPWR VGND _10251_ sg13g2_xnor2_1
X_17381_ _10249_ _10251_ VPWR VGND _10252_ sg13g2_nor2_1
X_17382_ _08568_ _10180_ _10181_ _10252_ VPWR VGND 
+ _10253_
+ sg13g2_a22oi_1
X_17383_ _10249_ _10251_ _08930_ VPWR VGND _10254_ sg13g2_a21oi_1
X_17384_ _10120_ _10147_ VPWR VGND _10255_ sg13g2_or2_1
X_17385_ _10255_ VPWR VGND _10256_ sg13g2_buf_1
X_17386_ _08463_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[13]\ VPWR VGND _10257_ sg13g2_xnor2_1
X_17387_ _10256_ _10257_ VPWR VGND _10258_ sg13g2_xnor2_1
X_17388_ _10181_ _10254_ _10258_ _08646_ VPWR VGND 
+ _10259_
+ sg13g2_a22oi_1
X_17389_ _10253_ _10259_ VPWR VGND _10260_ sg13g2_nand2_1
X_17390_ _08849_ _10148_ VPWR VGND _10261_ sg13g2_nor2_1
X_17391_ _08645_ _10256_ _10261_ VPWR VGND _10262_ sg13g2_o21ai_1
X_17392_ _10256_ _10257_ VPWR VGND _10263_ sg13g2_nor2_1
X_17393_ _10153_ _08676_ VPWR VGND _10264_ sg13g2_xnor2_1
X_17394_ _10263_ _10264_ VPWR VGND _10265_ sg13g2_nor2_1
X_17395_ _10147_ _10150_ _08645_ VPWR VGND _10266_ sg13g2_o21ai_1
X_17396_ _10149_ _10266_ _08843_ VPWR VGND _10267_ sg13g2_a21o_1
X_17397_ _08644_ _10149_ _10264_ VPWR VGND _10268_ sg13g2_o21ai_1
X_17398_ _10268_ VPWR VGND _10269_ sg13g2_inv_1
X_17399_ _10262_ _10265_ _10267_ _10269_ VPWR VGND 
+ _10270_
+ sg13g2_a22oi_1
X_17400_ _10173_ _10260_ _10270_ VPWR VGND _10271_ sg13g2_nand3_1
X_17401_ _08954_ _10260_ _10270_ VPWR VGND _10272_ sg13g2_nand3_1
X_17402_ _08954_ _10173_ VPWR VGND _10273_ sg13g2_nand2_1
X_17403_ _10177_ _10271_ _10272_ _10273_ VPWR VGND 
+ _10274_
+ sg13g2_nand4_1
X_17404_ _08729_ _10170_ _10171_ _10274_ VPWR VGND 
+ _10275_
+ sg13g2_a22oi_1
X_17405_ _10167_ _10168_ _10275_ VPWR VGND _10276_ sg13g2_a21oi_1
X_17406_ _08709_ _10166_ VPWR VGND _10277_ sg13g2_and2_1
X_17407_ _10164_ _10163_ _08740_ VPWR VGND _10278_ sg13g2_o21ai_1
X_17408_ _10164_ _10163_ VPWR VGND _10279_ sg13g2_nand2_1
X_17409_ _10278_ _10279_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2673_o\ VPWR VGND _10280_ sg13g2_a21oi_1
X_17410_ _08759_ _10280_ VPWR VGND _10281_ sg13g2_nor2_1
X_17411_ _10276_ _10277_ _10281_ VPWR VGND _10282_ sg13g2_o21ai_1
X_17412_ _10112_ VPWR VGND _10283_ sg13g2_inv_1
X_17413_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2671_o[0]\ VPWR VGND _10284_ sg13g2_buf_1
X_17414_ _07801_ VPWR VGND _10285_ sg13g2_buf_1
X_17415_ _10284_ _10285_ VPWR VGND _10286_ sg13g2_nand2_1
X_17416_ _10283_ _08977_ _10286_ VPWR VGND _10287_ sg13g2_o21ai_1
X_17417_ _10282_ _10287_ VPWR VGND _00509_ sg13g2_and2_1
X_17418_ _10115_ VPWR VGND _10288_ sg13g2_inv_1
X_17419_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2671_o[1]\ VPWR VGND _10289_ sg13g2_buf_1
X_17420_ _10289_ _10285_ VPWR VGND _10290_ sg13g2_nand2_1
X_17421_ _10288_ _08977_ _10290_ VPWR VGND _10291_ sg13g2_o21ai_1
X_17422_ _10282_ _10291_ VPWR VGND _00510_ sg13g2_and2_1
X_17423_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[17]\ VPWR VGND _10292_ sg13g2_buf_1
X_17424_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[16]\ VPWR VGND _10293_ sg13g2_buf_1
X_17425_ _08724_ _10293_ VPWR VGND _10294_ sg13g2_and2_1
X_17426_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[15]\ VPWR VGND _10295_ sg13g2_buf_1
X_17427_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[13]\ VPWR VGND _10296_ sg13g2_buf_1
X_17428_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[14]\ VPWR VGND _10297_ sg13g2_buf_1
X_17429_ _08650_ _10297_ VPWR VGND _10298_ sg13g2_nor2_1
X_17430_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[12]\ VPWR VGND _10299_ sg13g2_buf_1
X_17431_ _08609_ _10299_ VPWR VGND _10300_ sg13g2_nor2_1
X_17432_ _10298_ _10300_ VPWR VGND _10301_ sg13g2_nor2_1
X_17433_ _10296_ _10301_ VPWR VGND _10302_ sg13g2_nand2_1
X_17434_ _08660_ _10301_ VPWR VGND _10303_ sg13g2_nand2_1
X_17435_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[11]\ VPWR VGND _10304_ sg13g2_buf_1
X_17436_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[9]\ VPWR VGND _10305_ sg13g2_buf_1
X_17437_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[8]\ VPWR VGND _10306_ sg13g2_buf_1
X_17438_ _08417_ _10306_ VPWR VGND _10307_ sg13g2_or2_1
X_17439_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[6]\ VPWR VGND _10308_ sg13g2_buf_1
X_17440_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[7]\ VPWR VGND _10309_ sg13g2_buf_1
X_17441_ _08425_ _10308_ _10309_ VPWR VGND _10310_ sg13g2_a21oi_1
X_17442_ _08426_ _10309_ _10308_ VPWR VGND _10311_ sg13g2_nand3_1
X_17443_ _09361_ _10310_ _10311_ VPWR VGND _10312_ sg13g2_o21ai_1
X_17444_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[10]\ VPWR VGND _10313_ sg13g2_buf_1
X_17445_ _08433_ _10313_ _10306_ _08436_ VPWR VGND 
+ _10314_
+ sg13g2_a22oi_1
X_17446_ _10314_ VPWR VGND _10315_ sg13g2_inv_1
X_17447_ _08412_ _10305_ _10307_ _10312_ _10315_ VPWR 
+ VGND
+ _10316_ sg13g2_a221oi_1
X_17448_ _10316_ VPWR VGND _10317_ sg13g2_buf_1
X_17449_ _10305_ VPWR VGND _10318_ sg13g2_inv_1
X_17450_ _08434_ _10313_ VPWR VGND _10319_ sg13g2_nand2_1
X_17451_ _08443_ _10318_ _10319_ VPWR VGND _10320_ sg13g2_nand3_1
X_17452_ _08441_ _10313_ _10320_ VPWR VGND _10321_ sg13g2_o21ai_1
X_17453_ _10317_ _10321_ _08638_ VPWR VGND _10322_ sg13g2_o21ai_1
X_17454_ _08638_ _10317_ _10321_ VPWR VGND _10323_ sg13g2_nor3_1
X_17455_ _08455_ _10299_ _10304_ _10322_ _10323_ VPWR 
+ VGND
+ _10324_ sg13g2_a221oi_1
X_17456_ _10324_ VPWR VGND _10325_ sg13g2_buf_1
X_17457_ _10302_ _10303_ _10325_ VPWR VGND _10326_ sg13g2_a21oi_1
X_17458_ _10296_ VPWR VGND _10327_ sg13g2_inv_1
X_17459_ _08848_ _10327_ _10298_ VPWR VGND _10328_ sg13g2_nor3_1
X_17460_ _08652_ _10297_ _10328_ VPWR VGND _10329_ sg13g2_a21oi_1
X_17461_ _10326_ _10329_ VPWR VGND _10330_ sg13g2_nand2b_1
X_17462_ _10295_ _10330_ VPWR VGND _10331_ sg13g2_nor2_1
X_17463_ _10295_ _10330_ _08667_ VPWR VGND _10332_ sg13g2_a21oi_1
X_17464_ _10331_ _10332_ VPWR VGND _10333_ sg13g2_nor2_1
X_17465_ _10294_ _10333_ VPWR VGND _10334_ sg13g2_nor2_1
X_17466_ _09205_ _10293_ VPWR VGND _10335_ sg13g2_or2_1
X_17467_ _10334_ _10335_ VPWR VGND _10336_ sg13g2_nor2b_1
X_17468_ _10292_ _10336_ _08740_ VPWR VGND _10337_ sg13g2_o21ai_1
X_17469_ _10292_ _10336_ VPWR VGND _10338_ sg13g2_nand2_1
X_17470_ _10337_ _10338_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2676_o\ VPWR VGND _10339_ sg13g2_a21o_1
X_17471_ _10294_ _10333_ _10335_ VPWR VGND _10340_ sg13g2_o21ai_1
X_17472_ _08738_ _10292_ VPWR VGND _10341_ sg13g2_xnor2_1
X_17473_ _10340_ _10341_ VPWR VGND _10342_ sg13g2_xnor2_1
X_17474_ _08708_ _10342_ VPWR VGND _10343_ sg13g2_nand2_1
X_17475_ _08702_ _08728_ VPWR VGND _10344_ sg13g2_nor2_1
X_17476_ _08725_ _10293_ VPWR VGND _10345_ sg13g2_xor2_1
X_17477_ _10333_ _10345_ VPWR VGND _10346_ sg13g2_xnor2_1
X_17478_ _08702_ _10344_ _10346_ VPWR VGND _10347_ sg13g2_mux2_1
X_17479_ _08940_ _10295_ VPWR VGND _10348_ sg13g2_xnor2_1
X_17480_ _10330_ _10348_ VPWR VGND _10349_ sg13g2_xnor2_1
X_17481_ _08551_ _10306_ VPWR VGND _10350_ sg13g2_nor2_1
X_17482_ _08551_ _10306_ _10312_ VPWR VGND _10351_ sg13g2_a21oi_1
X_17483_ _10350_ _10351_ VPWR VGND _10352_ sg13g2_nor2_1
X_17484_ _10305_ _10352_ VPWR VGND _10353_ sg13g2_nand2_1
X_17485_ _10305_ _10352_ VPWR VGND _10354_ sg13g2_nor2_1
X_17486_ _08625_ _10353_ _10354_ VPWR VGND _10355_ sg13g2_a21oi_1
X_17487_ _08595_ _10313_ VPWR VGND _10356_ sg13g2_xor2_1
X_17488_ _10355_ _10356_ VPWR VGND _10357_ sg13g2_xnor2_1
X_17489_ _10313_ _08623_ VPWR VGND _10358_ sg13g2_xor2_1
X_17490_ _08577_ _10305_ _10352_ VPWR VGND _10359_ sg13g2_nor3_1
X_17491_ _08625_ _10354_ _10353_ _10044_ _10359_ VPWR 
+ VGND
+ _10360_ sg13g2_a221oi_1
X_17492_ _08861_ _10305_ VPWR VGND _10361_ sg13g2_nand2_1
X_17493_ _08577_ _10352_ _10361_ VPWR VGND _10362_ sg13g2_a21oi_1
X_17494_ _08584_ _10305_ VPWR VGND _10363_ sg13g2_xnor2_1
X_17495_ _10350_ _10351_ _10363_ VPWR VGND _10364_ sg13g2_nor3_1
X_17496_ _10362_ _10364_ _10358_ VPWR VGND _10365_ sg13g2_o21ai_1
X_17497_ _10358_ _10360_ _10365_ VPWR VGND _10366_ sg13g2_o21ai_1
X_17498_ _08469_ _10309_ VPWR VGND _10367_ sg13g2_xor2_1
X_17499_ _10367_ _08532_ VPWR VGND _10368_ sg13g2_nand2b_1
X_17500_ _10368_ VPWR VGND _10369_ sg13g2_buf_1
X_17501_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[252]\ VPWR VGND _10370_ sg13g2_buf_1
X_17502_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ VPWR VGND _10371_ sg13g2_buf_1
X_17503_ _10371_ _08882_ VPWR VGND _10372_ sg13g2_nand2b_1
X_17504_ _10370_ _10372_ VPWR VGND _10373_ sg13g2_nand2_1
X_17505_ _10370_ _10372_ _09061_ VPWR VGND _10374_ sg13g2_o21ai_1
X_17506_ _10373_ _10374_ VPWR VGND _10375_ sg13g2_nand2_1
X_17507_ _10308_ _10369_ _10375_ VPWR VGND _10376_ sg13g2_o21ai_1
X_17508_ _10308_ VPWR VGND _10377_ sg13g2_inv_1
X_17509_ _08556_ _10377_ VPWR VGND _10378_ sg13g2_nand2_1
X_17510_ _10369_ _10378_ _08543_ VPWR VGND _10379_ sg13g2_a21oi_1
X_17511_ _08534_ _10367_ _08557_ VPWR VGND _10380_ sg13g2_a21oi_1
X_17512_ _08516_ _10377_ _10380_ VPWR VGND _10381_ sg13g2_nor3_1
X_17513_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ VPWR VGND _10382_ sg13g2_inv_1
X_17514_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ VPWR VGND _10383_ sg13g2_buf_1
X_17515_ _08889_ _10383_ VPWR VGND _10384_ sg13g2_nor2_1
X_17516_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[248]\ VPWR VGND _10385_ sg13g2_buf_1
X_17517_ _10385_ _08891_ VPWR VGND _10386_ sg13g2_nand2b_1
X_17518_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ VPWR VGND _10387_ sg13g2_nor2b_1
X_17519_ _09071_ _10385_ VPWR VGND _10388_ sg13g2_nor2b_1
X_17520_ _08491_ _10383_ _10386_ _10387_ _10388_ VPWR 
+ VGND
+ _10389_ sg13g2_a221oi_1
X_17521_ _10384_ _10389_ VPWR VGND _10390_ sg13g2_or2_1
X_17522_ _10382_ _10390_ _08885_ VPWR VGND _10391_ sg13g2_o21ai_1
X_17523_ _10382_ _10390_ VPWR VGND _10392_ sg13g2_nand2_1
X_17524_ _08879_ _10370_ VPWR VGND _10393_ sg13g2_nor2b_1
X_17525_ _08884_ _10371_ _10391_ _10392_ _10393_ VPWR 
+ VGND
+ _10394_ sg13g2_a221oi_1
X_17526_ _10376_ _10379_ _10381_ _10394_ VPWR VGND 
+ _10395_
+ sg13g2_nor4_1
X_17527_ _08527_ _10367_ VPWR VGND _10396_ sg13g2_and2_1
X_17528_ _10306_ _10312_ VPWR VGND _10397_ sg13g2_xnor2_1
X_17529_ _09792_ _10397_ VPWR VGND _10398_ sg13g2_xor2_1
X_17530_ _10377_ _10396_ _10398_ VPWR VGND _10399_ sg13g2_a21oi_1
X_17531_ _08474_ _10308_ VPWR VGND _10400_ sg13g2_nand2_1
X_17532_ _10308_ _10192_ _10400_ VPWR VGND _10401_ sg13g2_o21ai_1
X_17533_ _10369_ _10401_ _10396_ VPWR VGND _10402_ sg13g2_a21o_1
X_17534_ _08508_ _10377_ _10369_ VPWR VGND _10403_ sg13g2_nand3_1
X_17535_ _10192_ _10367_ _08533_ VPWR VGND _10404_ sg13g2_a21oi_1
X_17536_ _10192_ _10367_ VPWR VGND _10405_ sg13g2_nor2_1
X_17537_ _10404_ _10405_ _10308_ VPWR VGND _10406_ sg13g2_o21ai_1
X_17538_ _08543_ _10403_ _10406_ VPWR VGND _10407_ sg13g2_nand3_1
X_17539_ _08543_ _10402_ _10407_ VPWR VGND _10408_ sg13g2_o21ai_1
X_17540_ _10399_ _10408_ VPWR VGND _10409_ sg13g2_nand2_1
X_17541_ _10352_ _10363_ VPWR VGND _10410_ sg13g2_xor2_1
X_17542_ _10124_ _10397_ VPWR VGND _10411_ sg13g2_xnor2_1
X_17543_ _08921_ _10410_ _10411_ _08605_ VPWR VGND 
+ _10412_
+ sg13g2_a22oi_1
X_17544_ _10395_ _10409_ _10412_ VPWR VGND _10413_ sg13g2_o21ai_1
X_17545_ _09048_ _10357_ _10366_ _10413_ VPWR VGND 
+ _10414_
+ sg13g2_a22oi_1
X_17546_ _10317_ _10321_ VPWR VGND _10415_ sg13g2_nor2_1
X_17547_ _08617_ _10304_ VPWR VGND _10416_ sg13g2_xnor2_1
X_17548_ _10415_ _10416_ VPWR VGND _10417_ sg13g2_xnor2_1
X_17549_ _10304_ _10322_ _10323_ VPWR VGND _10418_ sg13g2_a21oi_1
X_17550_ _08570_ _10299_ VPWR VGND _10419_ sg13g2_xnor2_1
X_17551_ _10418_ _10419_ VPWR VGND _10420_ sg13g2_xnor2_1
X_17552_ _09106_ _10420_ VPWR VGND _10421_ sg13g2_xnor2_1
X_17553_ _10414_ _10417_ _10421_ VPWR VGND _10422_ sg13g2_a21oi_1
X_17554_ _10414_ _10417_ _08930_ VPWR VGND _10423_ sg13g2_o21ai_1
X_17555_ _10325_ _10300_ _10327_ VPWR VGND _10424_ sg13g2_o21ai_1
X_17556_ _10327_ _10325_ _10300_ VPWR VGND _10425_ sg13g2_nor3_1
X_17557_ _08463_ _10424_ _10425_ VPWR VGND _10426_ sg13g2_a21oi_1
X_17558_ _08653_ _10297_ VPWR VGND _10427_ sg13g2_xnor2_1
X_17559_ _10426_ _10427_ VPWR VGND _10428_ sg13g2_xnor2_1
X_17560_ _10325_ _10300_ VPWR VGND _10429_ sg13g2_nor2_1
X_17561_ _08463_ _10296_ VPWR VGND _10430_ sg13g2_xnor2_1
X_17562_ _10429_ _10430_ VPWR VGND _10431_ sg13g2_xnor2_1
X_17563_ _08568_ _10420_ VPWR VGND _10432_ sg13g2_nand2_1
X_17564_ _10431_ _10432_ VPWR VGND _10433_ sg13g2_nand2_1
X_17565_ _08684_ _10428_ _10433_ VPWR VGND _10434_ sg13g2_a21o_1
X_17566_ _08644_ _10432_ VPWR VGND _10435_ sg13g2_nand2_1
X_17567_ _08684_ _10428_ _10435_ VPWR VGND _10436_ sg13g2_a21o_1
X_17568_ _10422_ _10423_ _10434_ _10436_ VPWR VGND 
+ _10437_
+ sg13g2_a22oi_1
X_17569_ _09720_ _10428_ VPWR VGND _10438_ sg13g2_xnor2_1
X_17570_ _08844_ _10431_ VPWR VGND _10439_ sg13g2_nand2_1
X_17571_ _08684_ _10428_ _10438_ _10439_ VPWR VGND 
+ _10440_
+ sg13g2_a22oi_1
X_17572_ _10437_ _10440_ VPWR VGND _10441_ sg13g2_or2_1
X_17573_ _08681_ _10349_ _10441_ VPWR VGND _10442_ sg13g2_a21o_1
X_17574_ _08680_ _10349_ VPWR VGND _10443_ sg13g2_nor2_1
X_17575_ _08708_ _10342_ _10346_ _08728_ _10443_ VPWR 
+ VGND
+ _10444_ sg13g2_a221oi_1
X_17576_ _08741_ _08707_ VPWR VGND _10445_ sg13g2_nor2_1
X_17577_ _08742_ _10445_ _10342_ VPWR VGND _10446_ sg13g2_mux2_1
X_17578_ _10343_ _10347_ _10442_ _10444_ _10446_ VPWR 
+ VGND
+ _10447_ sg13g2_a221oi_1
X_17579_ _07932_ _10339_ _10447_ VPWR VGND _10448_ sg13g2_nand3_1
X_17580_ _10284_ VPWR VGND _10449_ sg13g2_inv_1
X_17581_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2674_o[0]\ VPWR VGND _10450_ sg13g2_buf_4
X_17582_ _10450_ _10285_ VPWR VGND _10451_ sg13g2_nand2_1
X_17583_ _10449_ _08977_ _10451_ VPWR VGND _10452_ sg13g2_o21ai_1
X_17584_ _10448_ _10452_ VPWR VGND _00511_ sg13g2_and2_1
X_17585_ _10289_ VPWR VGND _10453_ sg13g2_inv_1
X_17586_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2674_o[1]\ VPWR VGND _10454_ sg13g2_buf_1
X_17587_ _10454_ VPWR VGND _10455_ sg13g2_buf_4
X_17588_ _10455_ _10285_ VPWR VGND _10456_ sg13g2_nand2_1
X_17589_ _10453_ _08977_ _10456_ VPWR VGND _10457_ sg13g2_o21ai_1
X_17590_ _10448_ _10457_ VPWR VGND _00512_ sg13g2_and2_1
X_17591_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n3499_o\ VPWR VGND _10458_ sg13g2_buf_2
X_17592_ _10458_ VPWR VGND _10459_ sg13g2_inv_1
X_17593_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[15]\ VPWR VGND _10460_ sg13g2_inv_1
X_17594_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[13]\ VPWR VGND _10461_ sg13g2_buf_1
X_17595_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[14]\ VPWR VGND _10462_ sg13g2_buf_1
X_17596_ _08650_ _10462_ VPWR VGND _10463_ sg13g2_nor2_1
X_17597_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[12]\ VPWR VGND _10464_ sg13g2_buf_1
X_17598_ _08453_ _10464_ VPWR VGND _10465_ sg13g2_or2_1
X_17599_ _10465_ VPWR VGND _10466_ sg13g2_buf_1
X_17600_ _10463_ _10466_ VPWR VGND _10467_ sg13g2_nor2b_1
X_17601_ _10461_ _10467_ VPWR VGND _10468_ sg13g2_and2_1
X_17602_ _08461_ _10467_ VPWR VGND _10469_ sg13g2_and2_1
X_17603_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[9]\ VPWR VGND _10470_ sg13g2_buf_1
X_17604_ _10470_ VPWR VGND _10471_ sg13g2_inv_1
X_17605_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[8]\ VPWR VGND _10472_ sg13g2_inv_1
X_17606_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[6]\ VPWR VGND _10473_ sg13g2_buf_1
X_17607_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[7]\ VPWR VGND _10474_ sg13g2_buf_1
X_17608_ _08425_ _10473_ _10474_ VPWR VGND _10475_ sg13g2_a21o_1
X_17609_ _08425_ _10474_ _10473_ VPWR VGND _10476_ sg13g2_and3_1
X_17610_ _08416_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[8]\ _10475_ _08422_ _10476_ VPWR 
+ VGND
+ _10477_ sg13g2_a221oi_1
X_17611_ _08443_ _10471_ _10472_ _10124_ _10477_ VPWR 
+ VGND
+ _10478_ sg13g2_a221oi_1
X_17612_ _10478_ VPWR VGND _10479_ sg13g2_buf_1
X_17613_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[10]\ VPWR VGND _10480_ sg13g2_buf_1
X_17614_ _08434_ _10480_ VPWR VGND _10481_ sg13g2_nand2_1
X_17615_ _08443_ _10471_ _10481_ VPWR VGND _10482_ sg13g2_o21ai_1
X_17616_ _08433_ _10480_ VPWR VGND _10483_ sg13g2_or2_1
X_17617_ _10483_ VPWR VGND _10484_ sg13g2_buf_1
X_17618_ _08406_ _10484_ VPWR VGND _10485_ sg13g2_and2_1
X_17619_ _10479_ _10482_ _10485_ VPWR VGND _10486_ sg13g2_o21ai_1
X_17620_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[11]\ VPWR VGND _10487_ sg13g2_buf_1
X_17621_ _10487_ _10484_ VPWR VGND _10488_ sg13g2_and2_1
X_17622_ _10479_ _10482_ _10488_ VPWR VGND _10489_ sg13g2_o21ai_1
X_17623_ _08454_ _10464_ _10487_ _08406_ VPWR VGND 
+ _10490_
+ sg13g2_a22oi_1
X_17624_ _10486_ _10489_ _10490_ VPWR VGND _10491_ sg13g2_nand3_1
X_17625_ _10491_ VPWR VGND _10492_ sg13g2_buf_1
X_17626_ _10468_ _10469_ _10492_ VPWR VGND _10493_ sg13g2_o21ai_1
X_17627_ _10461_ VPWR VGND _10494_ sg13g2_inv_1
X_17628_ _08848_ _10494_ _10463_ VPWR VGND _10495_ sg13g2_nor3_1
X_17629_ _08652_ _10462_ _10495_ VPWR VGND _10496_ sg13g2_a21oi_1
X_17630_ _10460_ _10493_ _10496_ VPWR VGND _10497_ sg13g2_nand3_1
X_17631_ _10493_ _10496_ _10460_ VPWR VGND _10498_ sg13g2_a21oi_1
X_17632_ _08667_ _10497_ _10498_ VPWR VGND _10499_ sg13g2_a21o_1
X_17633_ _10499_ VPWR VGND _10500_ sg13g2_buf_1
X_17634_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[16]\ VPWR VGND _10501_ sg13g2_buf_1
X_17635_ _08701_ _10501_ VPWR VGND _10502_ sg13g2_and2_1
X_17636_ _08724_ _10501_ VPWR VGND _10503_ sg13g2_or2_1
X_17637_ _10502_ _10503_ VPWR VGND _10504_ sg13g2_nor2b_1
X_17638_ _10500_ _10504_ VPWR VGND _10505_ sg13g2_xnor2_1
X_17639_ _10501_ _08704_ VPWR VGND _10506_ sg13g2_xor2_1
X_17640_ _10500_ _10506_ VPWR VGND _10507_ sg13g2_xnor2_1
X_17641_ _10493_ _10496_ VPWR VGND _10508_ sg13g2_nand2_1
X_17642_ _08668_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[15]\ VPWR VGND _10509_ sg13g2_xnor2_1
X_17643_ _10508_ _10509_ VPWR VGND _10510_ sg13g2_xnor2_1
X_17644_ _08680_ _10510_ VPWR VGND _10511_ sg13g2_nand2_1
X_17645_ _09720_ _08683_ VPWR VGND _10512_ sg13g2_nor2_1
X_17646_ _10492_ _10466_ _10461_ VPWR VGND _10513_ sg13g2_a21oi_1
X_17647_ _10461_ _10492_ _10466_ VPWR VGND _10514_ sg13g2_nand3_1
X_17648_ _08849_ _10513_ _10514_ VPWR VGND _10515_ sg13g2_o21ai_1
X_17649_ _08653_ _10462_ VPWR VGND _10516_ sg13g2_xnor2_1
X_17650_ _10515_ _10516_ VPWR VGND _10517_ sg13g2_xnor2_1
X_17651_ _10512_ _09720_ _10517_ VPWR VGND _10518_ sg13g2_mux2_1
X_17652_ _08680_ _10510_ _10518_ VPWR VGND _10519_ sg13g2_o21ai_1
X_17653_ _10507_ _10511_ _10519_ VPWR VGND _10520_ sg13g2_nand3_1
X_17654_ _10510_ VPWR VGND _10521_ sg13g2_inv_1
X_17655_ _10492_ _10466_ VPWR VGND _10522_ sg13g2_nand2_1
X_17656_ _08843_ _10461_ VPWR VGND _10523_ sg13g2_xor2_1
X_17657_ _10522_ _10523_ VPWR VGND _10524_ sg13g2_xnor2_1
X_17658_ _10479_ _10482_ _10484_ VPWR VGND _10525_ sg13g2_o21ai_1
X_17659_ _10487_ _10525_ VPWR VGND _10526_ sg13g2_nor2b_1
X_17660_ _08639_ _10489_ _10526_ VPWR VGND _10527_ sg13g2_a21o_1
X_17661_ _10464_ _10527_ VPWR VGND _10528_ sg13g2_xor2_1
X_17662_ _10064_ _10063_ _10528_ VPWR VGND _10529_ sg13g2_mux2_1
X_17663_ _10517_ _08684_ VPWR VGND _10530_ sg13g2_nand2b_1
X_17664_ _10524_ _10529_ _10530_ VPWR VGND _10531_ sg13g2_nand3_1
X_17665_ _09229_ _10529_ _10530_ VPWR VGND _10532_ sg13g2_nand3_1
X_17666_ _08617_ _10487_ VPWR VGND _10533_ sg13g2_xor2_1
X_17667_ _10525_ _10533_ VPWR VGND _10534_ sg13g2_xnor2_1
X_17668_ _10124_ _10472_ _10477_ VPWR VGND _10535_ sg13g2_a21oi_1
X_17669_ _08590_ _10535_ _10470_ VPWR VGND _10536_ sg13g2_a21o_1
X_17670_ _08861_ _10535_ _10536_ VPWR VGND _10537_ sg13g2_o21ai_1
X_17671_ _08595_ _10480_ VPWR VGND _10538_ sg13g2_xnor2_1
X_17672_ _10537_ _10538_ VPWR VGND _10539_ sg13g2_xnor2_1
X_17673_ _09048_ _10539_ VPWR VGND _10540_ sg13g2_nand2_1
X_17674_ _10534_ _10540_ VPWR VGND _10541_ sg13g2_nand2_1
X_17675_ _08930_ _10540_ VPWR VGND _10542_ sg13g2_nand2_1
X_17676_ _00074_ _10539_ VPWR VGND _10543_ sg13g2_xor2_1
X_17677_ _10473_ VPWR VGND _10544_ sg13g2_inv_1
X_17678_ _08578_ _10474_ VPWR VGND _10545_ sg13g2_xor2_1
X_17679_ _08534_ _10545_ _08556_ VPWR VGND _10546_ sg13g2_a21oi_1
X_17680_ _08516_ _10544_ _10546_ VPWR VGND _10547_ sg13g2_nor3_1
X_17681_ _10545_ _08533_ VPWR VGND _10548_ sg13g2_nand2b_1
X_17682_ _10548_ VPWR VGND _10549_ sg13g2_buf_1
X_17683_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _08879_ VPWR VGND _10550_ sg13g2_nand2b_1
X_17684_ _10473_ _10549_ _10550_ VPWR VGND _10551_ sg13g2_o21ai_1
X_17685_ _08557_ _10544_ VPWR VGND _10552_ sg13g2_nand2_1
X_17686_ _10549_ _10552_ _08543_ VPWR VGND _10553_ sg13g2_a21oi_1
X_17687_ _10547_ _10551_ _10553_ VPWR VGND _10554_ sg13g2_nor3_1
X_17688_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ VPWR VGND _10555_ sg13g2_inv_1
X_17689_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ VPWR VGND _10556_ sg13g2_inv_1
X_17690_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ _08892_ VPWR VGND _10557_ sg13g2_nand2b_1
X_17691_ _08894_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ VPWR VGND _10558_ sg13g2_nor2b_1
X_17692_ _08892_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ VPWR VGND _10559_ sg13g2_nor2b_1
X_17693_ _08889_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ _10557_ _10558_ _10559_ VPWR 
+ VGND
+ _10560_ sg13g2_a221oi_1
X_17694_ _08885_ _10555_ _10556_ _08888_ _10560_ VPWR 
+ VGND
+ _10561_ sg13g2_a221oi_1
X_17695_ _08487_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _08884_ _10561_ VPWR 
+ VGND
+ _10562_ sg13g2_a221oi_1
X_17696_ _08884_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ VPWR VGND _10563_ sg13g2_nor2_1
X_17697_ _09061_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ VPWR VGND _10564_ sg13g2_nand2_1
X_17698_ _10562_ _10563_ _10564_ VPWR VGND _10565_ sg13g2_o21ai_1
X_17699_ _10554_ _10565_ VPWR VGND _10566_ sg13g2_nand2_1
X_17700_ _08872_ _10545_ VPWR VGND _10567_ sg13g2_and2_1
X_17701_ _08534_ _10192_ _10545_ VPWR VGND _10568_ sg13g2_a21oi_1
X_17702_ _10193_ _10568_ _10473_ VPWR VGND _10569_ sg13g2_o21ai_1
X_17703_ _08508_ _10544_ _10549_ VPWR VGND _10570_ sg13g2_nand3_1
X_17704_ _08543_ _10569_ _10570_ VPWR VGND _10571_ sg13g2_nand3_1
X_17705_ _08508_ _10473_ VPWR VGND _10572_ sg13g2_nand2_1
X_17706_ _10473_ _10192_ _10572_ VPWR VGND _10573_ sg13g2_o21ai_1
X_17707_ _10549_ _10573_ _10567_ VPWR VGND _10574_ sg13g2_a21oi_1
X_17708_ _08516_ _10574_ VPWR VGND _10575_ sg13g2_nand2_1
X_17709_ _08867_ _10475_ _10476_ VPWR VGND _10576_ sg13g2_a21oi_1
X_17710_ _08551_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[8]\ VPWR VGND _10577_ sg13g2_xnor2_1
X_17711_ _10576_ _10577_ VPWR VGND _10578_ sg13g2_xnor2_1
X_17712_ _08549_ _10578_ VPWR VGND _10579_ sg13g2_xor2_1
X_17713_ _10544_ _10567_ _10571_ _10575_ _10579_ VPWR 
+ VGND
+ _10580_ sg13g2_a221oi_1
X_17714_ _08861_ _10470_ VPWR VGND _10581_ sg13g2_xnor2_1
X_17715_ _10535_ _10581_ VPWR VGND _10582_ sg13g2_xnor2_1
X_17716_ _08605_ _10578_ VPWR VGND _10583_ sg13g2_nand2_1
X_17717_ _10582_ _10583_ VPWR VGND _10584_ sg13g2_nand2_1
X_17718_ _10566_ _10580_ _10584_ VPWR VGND _10585_ sg13g2_a21oi_1
X_17719_ _08605_ VPWR VGND _10586_ sg13g2_buf_1
X_17720_ _10586_ _10578_ _10580_ _10566_ _08921_ VPWR 
+ VGND
+ _10587_ sg13g2_a221oi_1
X_17721_ _08577_ _10582_ VPWR VGND _10588_ sg13g2_and2_1
X_17722_ _10543_ _10585_ _10587_ _10588_ VPWR VGND 
+ _10589_
+ sg13g2_nor4_1
X_17723_ _10541_ _10542_ _10589_ VPWR VGND _10590_ sg13g2_a21oi_1
X_17724_ _08612_ _10528_ VPWR VGND _10591_ sg13g2_xnor2_1
X_17725_ _08930_ _10534_ _10591_ VPWR VGND _10592_ sg13g2_a21oi_1
X_17726_ _10590_ _10592_ VPWR VGND _10593_ sg13g2_nor2b_1
X_17727_ _08955_ _10521_ _10531_ _10532_ _10593_ VPWR 
+ VGND
+ _10594_ sg13g2_a221oi_1
X_17728_ _09229_ _10524_ _10530_ VPWR VGND _10595_ sg13g2_nand3_1
X_17729_ _08955_ _10521_ _10595_ VPWR VGND _10596_ sg13g2_a21oi_1
X_17730_ _10520_ _10594_ _10596_ VPWR VGND _10597_ sg13g2_nor3_1
X_17731_ _08729_ _10505_ _10597_ VPWR VGND _10598_ sg13g2_a21oi_1
X_17732_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3011_o\ VPWR VGND _10599_ sg13g2_buf_1
X_17733_ _10599_ _08758_ _08745_ VPWR VGND _10600_ sg13g2_o21ai_1
X_17734_ _08740_ _08741_ _10600_ VPWR VGND _10601_ sg13g2_o21ai_1
X_17735_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[17]\ VPWR VGND _10602_ sg13g2_buf_1
X_17736_ _10500_ _10502_ _10503_ VPWR VGND _10603_ sg13g2_o21ai_1
X_17737_ _10603_ VPWR VGND _10604_ sg13g2_buf_1
X_17738_ _10602_ _10604_ VPWR VGND _10605_ sg13g2_xnor2_1
X_17739_ _10599_ _08758_ _10602_ VPWR VGND _10606_ sg13g2_o21ai_1
X_17740_ _10602_ VPWR VGND _10607_ sg13g2_inv_1
X_17741_ _10607_ _10604_ VPWR VGND _10608_ sg13g2_nand2_1
X_17742_ _10604_ _10606_ _10608_ VPWR VGND _10609_ sg13g2_o21ai_1
X_17743_ _10601_ _10605_ _10609_ _08750_ VPWR VGND 
+ _10610_
+ sg13g2_a22oi_1
X_17744_ _08739_ _10602_ _10599_ _10604_ VPWR VGND 
+ _10611_
+ sg13g2_and4_1
X_17745_ _08822_ _10608_ VPWR VGND _10612_ sg13g2_nor2_1
X_17746_ _08739_ _10607_ _10599_ VPWR VGND _10613_ sg13g2_nand3_1
X_17747_ _08712_ _10602_ _10599_ VPWR VGND _10614_ sg13g2_nand3_1
X_17748_ _10613_ _10614_ _10604_ VPWR VGND _10615_ sg13g2_a21oi_1
X_17749_ _10611_ _10612_ _10615_ VPWR VGND _10616_ sg13g2_or3_1
X_17750_ _08709_ _10616_ _08759_ VPWR VGND _10617_ sg13g2_a21oi_1
X_17751_ _10598_ _10610_ _10617_ VPWR VGND _10618_ sg13g2_o21ai_1
X_17752_ _08759_ VPWR VGND _10619_ sg13g2_buf_1
X_17753_ _10450_ _10619_ VPWR VGND _10620_ sg13g2_nand2_1
X_17754_ _10459_ _10618_ _10620_ VPWR VGND _00513_ sg13g2_o21ai_1
X_17755_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n3496_o\ VPWR VGND _10621_ sg13g2_buf_1
X_17756_ _10621_ VPWR VGND _10622_ sg13g2_inv_1
X_17757_ _10455_ _10619_ VPWR VGND _10623_ sg13g2_nand2_1
X_17758_ _10622_ _10618_ _10623_ VPWR VGND _00514_ sg13g2_o21ai_1
X_17759_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2638_o[0]\ VPWR VGND _10624_ sg13g2_buf_1
X_17760_ _10624_ VPWR VGND _10625_ sg13g2_inv_1
X_17761_ _10625_ _08759_ VPWR VGND _10626_ sg13g2_nor2_1
X_17762_ _08403_ _08981_ _10626_ VPWR VGND _10627_ sg13g2_a21oi_1
X_17763_ _08758_ VPWR VGND _10628_ sg13g2_buf_1
X_17764_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2640_o\ VPWR VGND _10629_ sg13g2_buf_1
X_17765_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[17]\ VPWR VGND _10630_ sg13g2_inv_1
X_17766_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[15]\ VPWR VGND _10631_ sg13g2_buf_1
X_17767_ _10631_ VPWR VGND _10632_ sg13g2_inv_1
X_17768_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[16]\ VPWR VGND _10633_ sg13g2_buf_1
X_17769_ _10633_ VPWR VGND _10634_ sg13g2_inv_1
X_17770_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[13]\ VPWR VGND _10635_ sg13g2_buf_1
X_17771_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[12]\ VPWR VGND _10636_ sg13g2_buf_1
X_17772_ _08453_ _10636_ VPWR VGND _10637_ sg13g2_nor2_1
X_17773_ _10637_ VPWR VGND _10638_ sg13g2_inv_1
X_17774_ _10635_ _10638_ VPWR VGND _10639_ sg13g2_nor2_1
X_17775_ _08453_ _10636_ VPWR VGND _10640_ sg13g2_and2_1
X_17776_ _10640_ VPWR VGND _10641_ sg13g2_buf_1
X_17777_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[9]\ VPWR VGND _10642_ sg13g2_buf_1
X_17778_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[8]\ VPWR VGND _10643_ sg13g2_buf_1
X_17779_ _08415_ _10643_ VPWR VGND _10644_ sg13g2_or2_1
X_17780_ _10644_ VPWR VGND _10645_ sg13g2_buf_1
X_17781_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[6]\ VPWR VGND _10646_ sg13g2_buf_1
X_17782_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[7]\ VPWR VGND _10647_ sg13g2_buf_1
X_17783_ _08424_ _10646_ _10647_ VPWR VGND _10648_ sg13g2_a21oi_1
X_17784_ _08424_ _10647_ _10646_ VPWR VGND _10649_ sg13g2_nand3_1
X_17785_ _09361_ _10648_ _10649_ VPWR VGND _10650_ sg13g2_o21ai_1
X_17786_ _10650_ VPWR VGND _10651_ sg13g2_buf_1
X_17787_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[10]\ VPWR VGND _10652_ sg13g2_buf_1
X_17788_ _08415_ _10643_ VPWR VGND _10653_ sg13g2_and2_1
X_17789_ _10653_ VPWR VGND _10654_ sg13g2_buf_1
X_17790_ _08432_ _10652_ _10654_ VPWR VGND _10655_ sg13g2_a21o_1
X_17791_ _08412_ _10642_ _10645_ _10651_ _10655_ VPWR 
+ VGND
+ _10656_ sg13g2_a221oi_1
X_17792_ _10656_ VPWR VGND _10657_ sg13g2_buf_1
X_17793_ _08432_ _10652_ VPWR VGND _10658_ sg13g2_or2_1
X_17794_ _10658_ VPWR VGND _10659_ sg13g2_buf_1
X_17795_ _08433_ _10652_ VPWR VGND _10660_ sg13g2_nand2_1
X_17796_ _08412_ _10642_ VPWR VGND _10661_ sg13g2_nor2_1
X_17797_ _10660_ _10661_ VPWR VGND _10662_ sg13g2_nand2_1
X_17798_ _10659_ _10662_ VPWR VGND _10663_ sg13g2_nand2_1
X_17799_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[11]\ VPWR VGND _10664_ sg13g2_inv_1
X_17800_ _10657_ _10663_ _10664_ VPWR VGND _10665_ sg13g2_o21ai_1
X_17801_ _10635_ _10641_ _10665_ VPWR VGND _10666_ sg13g2_nor3_1
X_17802_ _10664_ _10657_ _10663_ VPWR VGND _10667_ sg13g2_nor3_1
X_17803_ _08407_ _10635_ _10641_ _10667_ VPWR VGND 
+ _10668_
+ sg13g2_nor4_1
X_17804_ _10639_ _10666_ _10668_ VPWR VGND _10669_ sg13g2_or3_1
X_17805_ _10669_ VPWR VGND _10670_ sg13g2_buf_1
X_17806_ _10641_ _10665_ VPWR VGND _10671_ sg13g2_or2_1
X_17807_ _08994_ _10641_ _10667_ VPWR VGND _10672_ sg13g2_or3_1
X_17808_ _10635_ _10638_ _10671_ _10672_ VPWR VGND 
+ _10673_
+ sg13g2_nand4_1
X_17809_ _08849_ _10670_ _10673_ VPWR VGND _10674_ sg13g2_o21ai_1
X_17810_ _10674_ VPWR VGND _10675_ sg13g2_buf_1
X_17811_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[14]\ VPWR VGND _10676_ sg13g2_buf_1
X_17812_ _08653_ _10676_ VPWR VGND _10677_ sg13g2_and2_1
X_17813_ _08653_ _10676_ VPWR VGND _10678_ sg13g2_or2_1
X_17814_ _10675_ _10677_ _10678_ VPWR VGND _10679_ sg13g2_o21ai_1
X_17815_ _10679_ VPWR VGND _10680_ sg13g2_buf_1
X_17816_ _08696_ _10632_ _10634_ _08716_ _10680_ VPWR 
+ VGND
+ _10681_ sg13g2_a221oi_1
X_17817_ _09205_ _10633_ VPWR VGND _10682_ sg13g2_nand2_1
X_17818_ _08669_ _10631_ _10633_ VPWR VGND _10683_ sg13g2_nand3_1
X_17819_ _08668_ _09205_ _10631_ VPWR VGND _10684_ sg13g2_nand3_1
X_17820_ _10682_ _10683_ _10684_ VPWR VGND _10685_ sg13g2_nand3_1
X_17821_ _10681_ _10685_ VPWR VGND _10686_ sg13g2_nor2_1
X_17822_ _10630_ _10686_ VPWR VGND _10687_ sg13g2_nor2_1
X_17823_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[17]\ _10681_ _10685_ VPWR VGND _10688_ sg13g2_nor3_1
X_17824_ _10629_ _10687_ _10688_ VPWR VGND _10689_ sg13g2_a21o_1
X_17825_ _10688_ _10687_ VPWR VGND _10690_ sg13g2_nor2_1
X_17826_ _10629_ _08745_ VPWR VGND _10691_ sg13g2_nand2_1
X_17827_ _08740_ _08742_ _10691_ VPWR VGND _10692_ sg13g2_o21ai_1
X_17828_ _08750_ _10689_ _10690_ _10692_ VPWR VGND 
+ _10693_
+ sg13g2_a22oi_1
X_17829_ _10632_ _10680_ VPWR VGND _10694_ sg13g2_nand2_1
X_17830_ _10632_ _10680_ _08696_ VPWR VGND _10695_ sg13g2_o21ai_1
X_17831_ _10694_ _10695_ VPWR VGND _10696_ sg13g2_nand2_1
X_17832_ _08725_ _10633_ VPWR VGND _10697_ sg13g2_xnor2_1
X_17833_ _10696_ _10697_ VPWR VGND _10698_ sg13g2_xnor2_1
X_17834_ _08702_ _10698_ VPWR VGND _10699_ sg13g2_xnor2_1
X_17835_ _08682_ _10676_ VPWR VGND _10700_ sg13g2_xor2_1
X_17836_ _10675_ _10700_ VPWR VGND _10701_ sg13g2_xnor2_1
X_17837_ _10657_ _10663_ VPWR VGND _10702_ sg13g2_nor2_1
X_17838_ _08408_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[11]\ VPWR VGND _10703_ sg13g2_xnor2_1
X_17839_ _10702_ _10703_ VPWR VGND _10704_ sg13g2_xor2_1
X_17840_ _08616_ _10667_ _10665_ VPWR VGND _10705_ sg13g2_o21ai_1
X_17841_ _08456_ _10636_ VPWR VGND _10706_ sg13g2_xnor2_1
X_17842_ _10705_ _10706_ VPWR VGND _10707_ sg13g2_xnor2_1
X_17843_ _08582_ _10642_ _10645_ _10651_ _10654_ VPWR 
+ VGND
+ _10708_ sg13g2_a221oi_1
X_17844_ _08589_ _10659_ _10660_ VPWR VGND _10709_ sg13g2_nand3_1
X_17845_ _10661_ _10708_ _10709_ VPWR VGND _10710_ sg13g2_nor3_1
X_17846_ _10659_ _10660_ _08860_ VPWR VGND _10711_ sg13g2_a21oi_1
X_17847_ _10661_ _10708_ _10711_ VPWR VGND _10712_ sg13g2_o21ai_1
X_17848_ _10710_ _10712_ VPWR VGND _10713_ sg13g2_nor2b_1
X_17849_ _08550_ _10643_ VPWR VGND _10714_ sg13g2_xor2_1
X_17850_ _10651_ _10714_ VPWR VGND _10715_ sg13g2_xnor2_1
X_17851_ _10645_ _10651_ _10654_ VPWR VGND _10716_ sg13g2_a21o_1
X_17852_ _10716_ VPWR VGND _10717_ sg13g2_buf_1
X_17853_ _08583_ _10642_ VPWR VGND _10718_ sg13g2_xor2_1
X_17854_ _10717_ _10718_ VPWR VGND _10719_ sg13g2_xnor2_1
X_17855_ _08604_ _10715_ _10719_ _08920_ VPWR VGND 
+ _10720_
+ sg13g2_a22oi_1
X_17856_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[22]\ VPWR VGND _10721_ sg13g2_inv_1
X_17857_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ VPWR VGND _10722_ sg13g2_inv_1
X_17858_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[20]\ VPWR VGND _10723_ sg13g2_buf_1
X_17859_ _10723_ _09071_ VPWR VGND _10724_ sg13g2_nand2b_1
X_17860_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ VPWR VGND _10725_ sg13g2_nor2b_1
X_17861_ _09071_ _10723_ VPWR VGND _10726_ sg13g2_nor2b_1
X_17862_ _08491_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ _10724_ _10725_ _10726_ VPWR 
+ VGND
+ _10727_ sg13g2_a221oi_1
X_17863_ _08485_ _10721_ _10722_ _08888_ _10727_ VPWR 
+ VGND
+ _10728_ sg13g2_a221oi_1
X_17864_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ VPWR VGND _10729_ sg13g2_buf_1
X_17865_ _08482_ _10729_ VPWR VGND _10730_ sg13g2_nand2_1
X_17866_ _08885_ _10721_ _10730_ VPWR VGND _10731_ sg13g2_o21ai_1
X_17867_ _08513_ _10646_ VPWR VGND _10732_ sg13g2_nand2_1
X_17868_ _08578_ _10647_ VPWR VGND _10733_ sg13g2_xnor2_1
X_17869_ _10732_ _10733_ VPWR VGND _10734_ sg13g2_xnor2_1
X_17870_ _08513_ _10646_ VPWR VGND _10735_ sg13g2_xnor2_1
X_17871_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[24]\ VPWR VGND _10736_ sg13g2_buf_1
X_17872_ _10729_ _08882_ VPWR VGND _10737_ sg13g2_nand2b_1
X_17873_ _08477_ _10736_ _10737_ VPWR VGND _10738_ sg13g2_o21ai_1
X_17874_ _08533_ _10734_ _10735_ _08556_ _10738_ VPWR 
+ VGND
+ _10739_ sg13g2_a221oi_1
X_17875_ _10728_ _10731_ _10739_ VPWR VGND _10740_ sg13g2_o21ai_1
X_17876_ _08548_ _10715_ VPWR VGND _10741_ sg13g2_xnor2_1
X_17877_ _08477_ _10736_ VPWR VGND _10742_ sg13g2_nand2_1
X_17878_ _10646_ _08901_ VPWR VGND _10743_ sg13g2_xnor2_1
X_17879_ _08556_ _10735_ VPWR VGND _10744_ sg13g2_and2_1
X_17880_ _08533_ _10734_ _10742_ _10743_ _10744_ VPWR 
+ VGND
+ _10745_ sg13g2_a221oi_1
X_17881_ _08534_ _10734_ VPWR VGND _10746_ sg13g2_nor2_1
X_17882_ _10745_ _10746_ VPWR VGND _10747_ sg13g2_nor2_1
X_17883_ _10740_ _10741_ _10747_ VPWR VGND _10748_ sg13g2_nand3_1
X_17884_ _10713_ _10720_ _10748_ VPWR VGND _10749_ sg13g2_nand3_1
X_17885_ _10702_ _10703_ VPWR VGND _10750_ sg13g2_xnor2_1
X_17886_ _08584_ _10642_ VPWR VGND _10751_ sg13g2_nand2_1
X_17887_ _08576_ _10717_ _10751_ VPWR VGND _10752_ sg13g2_a21oi_1
X_17888_ _10652_ _08622_ VPWR VGND _10753_ sg13g2_xnor2_1
X_17889_ _10717_ _10718_ _10753_ VPWR VGND _10754_ sg13g2_a21o_1
X_17890_ _08582_ _10642_ VPWR VGND _10755_ sg13g2_or2_1
X_17891_ _08574_ _10642_ VPWR VGND _10756_ sg13g2_or2_1
X_17892_ _10645_ _10651_ _10755_ _10756_ _10654_ VPWR 
+ VGND
+ _10757_ sg13g2_a221oi_1
X_17893_ _10654_ _10044_ VPWR VGND _10758_ sg13g2_nand2b_1
X_17894_ _10645_ _10651_ _10758_ VPWR VGND _10759_ sg13g2_a21oi_1
X_17895_ _08582_ _08575_ _10642_ VPWR VGND _10760_ sg13g2_nor3_1
X_17896_ _10760_ _10753_ VPWR VGND _10761_ sg13g2_nand2b_1
X_17897_ _10757_ _10759_ _10761_ VPWR VGND _10762_ sg13g2_or3_1
X_17898_ _10752_ _10754_ _10762_ VPWR VGND _10763_ sg13g2_o21ai_1
X_17899_ _08601_ _10750_ _10713_ _10763_ VPWR VGND 
+ _10764_
+ sg13g2_a22oi_1
X_17900_ _10749_ _10764_ VPWR VGND _10765_ sg13g2_and2_1
X_17901_ _08635_ _10704_ _10707_ _08568_ _10765_ VPWR 
+ VGND
+ _10766_ sg13g2_a221oi_1
X_17902_ _09106_ _08569_ VPWR VGND _10767_ sg13g2_nand2_1
X_17903_ _10767_ _10707_ VPWR VGND _10768_ sg13g2_nand2b_1
X_17904_ _09106_ _10707_ _10768_ VPWR VGND _10769_ sg13g2_o21ai_1
X_17905_ _10766_ _10769_ _08844_ VPWR VGND _10770_ sg13g2_o21ai_1
X_17906_ _10676_ _08840_ VPWR VGND _10771_ sg13g2_xnor2_1
X_17907_ _08849_ _10670_ VPWR VGND _10772_ sg13g2_nand2_1
X_17908_ _08849_ _10673_ VPWR VGND _10773_ sg13g2_nand2_1
X_17909_ _10635_ _10638_ _10671_ _10672_ VPWR VGND 
+ _10774_
+ sg13g2_and4_1
X_17910_ _10670_ _10774_ _08464_ VPWR VGND _10775_ sg13g2_o21ai_1
X_17911_ _10773_ _10771_ _10775_ VPWR VGND _10776_ sg13g2_nand3_1
X_17912_ _10771_ _10772_ _10776_ VPWR VGND _10777_ sg13g2_o21ai_1
X_17913_ _08464_ _10635_ VPWR VGND _10778_ sg13g2_nand2_1
X_17914_ _10675_ _10778_ _10771_ VPWR VGND _10779_ sg13g2_mux2_1
X_17915_ _08844_ _10766_ _10769_ _10779_ VPWR VGND 
+ _10780_
+ sg13g2_nor4_1
X_17916_ _08684_ _10701_ _10770_ _10777_ _10780_ VPWR 
+ VGND
+ _10781_ sg13g2_a221oi_1
X_17917_ _08940_ _10631_ VPWR VGND _10782_ sg13g2_xor2_1
X_17918_ _10680_ _10782_ VPWR VGND _10783_ sg13g2_xnor2_1
X_17919_ _08680_ _10781_ _10783_ VPWR VGND _10784_ sg13g2_a21o_1
X_17920_ _08681_ _10781_ _10784_ VPWR VGND _10785_ sg13g2_o21ai_1
X_17921_ _08729_ _10698_ _10699_ _10785_ VPWR VGND 
+ _10786_
+ sg13g2_a22oi_1
X_17922_ _10628_ _10693_ _10786_ VPWR VGND _10787_ sg13g2_nor3_1
X_17923_ _08740_ _10629_ _10690_ VPWR VGND _10788_ sg13g2_nand3_1
X_17924_ _10629_ VPWR VGND _10789_ sg13g2_inv_1
X_17925_ _08740_ _10789_ VPWR VGND _10790_ sg13g2_nor2_1
X_17926_ _08712_ _10688_ _10687_ _10790_ VPWR VGND 
+ _10791_
+ sg13g2_a22oi_1
X_17927_ _08709_ _07931_ VPWR VGND _10792_ sg13g2_nand2_1
X_17928_ _10788_ _10791_ _10792_ VPWR VGND _10793_ sg13g2_a21oi_1
X_17929_ _10627_ _10787_ _10793_ VPWR VGND _00515_ sg13g2_nor3_1
X_17930_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2638_o[1]\ VPWR VGND _10794_ sg13g2_buf_1
X_17931_ _10794_ VPWR VGND _10795_ sg13g2_inv_1
X_17932_ _10795_ _09710_ _08970_ VPWR VGND _10796_ sg13g2_mux2_1
X_17933_ _10787_ _10793_ _10796_ VPWR VGND _00516_ sg13g2_nor3_1
X_17934_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[16]\ VPWR VGND _10797_ sg13g2_buf_1
X_17935_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[15]\ VPWR VGND _10798_ sg13g2_buf_1
X_17936_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[11]\ VPWR VGND _10799_ sg13g2_buf_1
X_17937_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[12]\ VPWR VGND _10800_ sg13g2_buf_1
X_17938_ _08453_ _10800_ VPWR VGND _10801_ sg13g2_nor2_1
X_17939_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[10]\ VPWR VGND _10802_ sg13g2_buf_1
X_17940_ _08594_ _10802_ VPWR VGND _10803_ sg13g2_nor2_1
X_17941_ _10801_ _10803_ VPWR VGND _10804_ sg13g2_nor2_1
X_17942_ _10799_ _10804_ VPWR VGND _10805_ sg13g2_nand2_1
X_17943_ _08994_ _10804_ VPWR VGND _10806_ sg13g2_nand2_1
X_17944_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[8]\ VPWR VGND _10807_ sg13g2_buf_1
X_17945_ _08436_ _10807_ VPWR VGND _10808_ sg13g2_nor2_1
X_17946_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[6]\ VPWR VGND _10809_ sg13g2_buf_1
X_17947_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[7]\ VPWR VGND _10810_ sg13g2_buf_1
X_17948_ _08426_ _10809_ _10810_ VPWR VGND _10811_ sg13g2_a21o_1
X_17949_ _08426_ _10810_ _10809_ VPWR VGND _10812_ sg13g2_and3_1
X_17950_ _08417_ _10807_ _10811_ _08422_ _10812_ VPWR 
+ VGND
+ _10813_ sg13g2_a221oi_1
X_17951_ _10813_ VPWR VGND _10814_ sg13g2_buf_1
X_17952_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[9]\ VPWR VGND _10815_ sg13g2_buf_1
X_17953_ _10815_ VPWR VGND _10816_ sg13g2_inv_1
X_17954_ _10808_ _10814_ _10816_ VPWR VGND _10817_ sg13g2_o21ai_1
X_17955_ _10816_ _10808_ _10814_ VPWR VGND _10818_ sg13g2_nor3_1
X_17956_ _08582_ _10817_ _10818_ VPWR VGND _10819_ sg13g2_a21oi_1
X_17957_ _10805_ _10806_ _10819_ VPWR VGND _10820_ sg13g2_a21oi_1
X_17958_ _08406_ _10799_ VPWR VGND _10821_ sg13g2_nand2_1
X_17959_ _08441_ _10802_ VPWR VGND _10822_ sg13g2_nand2_1
X_17960_ _10801_ _10822_ VPWR VGND _10823_ sg13g2_nor2_1
X_17961_ _08407_ _10799_ _10823_ VPWR VGND _10824_ sg13g2_o21ai_1
X_17962_ _10801_ _10821_ _10824_ VPWR VGND _10825_ sg13g2_o21ai_1
X_17963_ _10825_ VPWR VGND _10826_ sg13g2_buf_1
X_17964_ _08609_ _10800_ VPWR VGND _10827_ sg13g2_and2_1
X_17965_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[14]\ VPWR VGND _10828_ sg13g2_buf_1
X_17966_ _08651_ _10828_ VPWR VGND _10829_ sg13g2_nand2_1
X_17967_ _10827_ _10829_ VPWR VGND _10830_ sg13g2_nand2b_1
X_17968_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[13]\ _10820_ _10826_ _10830_ VPWR VGND 
+ _10831_
+ sg13g2_nor4_1
X_17969_ _08660_ _10820_ _10826_ _10830_ VPWR VGND 
+ _10832_
+ sg13g2_nor4_1
X_17970_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[13]\ VPWR VGND _10833_ sg13g2_inv_1
X_17971_ _08848_ _10833_ _10829_ VPWR VGND _10834_ sg13g2_nand3_1
X_17972_ _08652_ _10828_ _10834_ VPWR VGND _10835_ sg13g2_o21ai_1
X_17973_ _10831_ _10832_ _10835_ VPWR VGND _10836_ sg13g2_nor3_1
X_17974_ _10798_ _10836_ _08667_ VPWR VGND _10837_ sg13g2_a21oi_1
X_17975_ _10798_ _10836_ VPWR VGND _10838_ sg13g2_nor2_1
X_17976_ _10837_ _10838_ VPWR VGND _10839_ sg13g2_nor2_1
X_17977_ _10797_ _10839_ VPWR VGND _10840_ sg13g2_xnor2_1
X_17978_ _08704_ _10840_ VPWR VGND _10841_ sg13g2_xnor2_1
X_17979_ _10820_ _10826_ _10827_ VPWR VGND _10842_ sg13g2_nor3_1
X_17980_ _08843_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[13]\ VPWR VGND _10843_ sg13g2_xor2_1
X_17981_ _10842_ _10843_ VPWR VGND _10844_ sg13g2_xnor2_1
X_17982_ _10819_ _10803_ _10822_ VPWR VGND _10845_ sg13g2_o21ai_1
X_17983_ _10845_ VPWR VGND _10846_ sg13g2_buf_1
X_17984_ _10799_ _10846_ VPWR VGND _10847_ sg13g2_nor2_1
X_17985_ _10799_ _10846_ VPWR VGND _10848_ sg13g2_nand2_1
X_17986_ _08639_ _10847_ _10848_ VPWR VGND _10849_ sg13g2_o21ai_1
X_17987_ _08570_ _10800_ VPWR VGND _10850_ sg13g2_xnor2_1
X_17988_ _10849_ _10850_ VPWR VGND _10851_ sg13g2_xnor2_1
X_17989_ _08569_ _10851_ VPWR VGND _10852_ sg13g2_nor2_1
X_17990_ _10800_ _08612_ VPWR VGND _10853_ sg13g2_xnor2_1
X_17991_ _10799_ _10846_ _08601_ VPWR VGND _10854_ sg13g2_a21oi_1
X_17992_ _10847_ _10854_ VPWR VGND _10855_ sg13g2_or2_1
X_17993_ _08635_ _10847_ _10855_ _08639_ VPWR VGND 
+ _10856_
+ sg13g2_a22oi_1
X_17994_ _08616_ _10799_ VPWR VGND _10857_ sg13g2_xor2_1
X_17995_ _10846_ _10857_ _10853_ VPWR VGND _10858_ sg13g2_a21oi_1
X_17996_ _08615_ _10846_ _10821_ VPWR VGND _10859_ sg13g2_a21o_1
X_17997_ _10846_ _10857_ VPWR VGND _10860_ sg13g2_xnor2_1
X_17998_ _10808_ _10814_ VPWR VGND _10861_ sg13g2_nor2_1
X_17999_ _08584_ _10815_ VPWR VGND _10862_ sg13g2_xor2_1
X_18000_ _08590_ _10815_ VPWR VGND _10863_ sg13g2_nand2_1
X_18001_ _08626_ _10861_ _10863_ VPWR VGND _10864_ sg13g2_a21oi_1
X_18002_ _10861_ _10862_ _10864_ VPWR VGND _10865_ sg13g2_a21oi_1
X_18003_ _10802_ _08623_ VPWR VGND _10866_ sg13g2_xor2_1
X_18004_ _10815_ _10861_ VPWR VGND _10867_ sg13g2_nor2_1
X_18005_ _08626_ _10818_ _10817_ VPWR VGND _10868_ sg13g2_o21ai_1
X_18006_ _08921_ _10867_ _10868_ _08625_ _10866_ VPWR 
+ VGND
+ _10869_ sg13g2_a221oi_1
X_18007_ _10865_ _10866_ _10869_ VPWR VGND _10870_ sg13g2_a21oi_1
X_18008_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[42]\ VPWR VGND _10871_ sg13g2_buf_1
X_18009_ _08884_ _10871_ VPWR VGND _10872_ sg13g2_nand2_1
X_18010_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ VPWR VGND _10873_ sg13g2_inv_1
X_18011_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[40]\ VPWR VGND _10874_ sg13g2_buf_1
X_18012_ _08889_ _10874_ VPWR VGND _10875_ sg13g2_nor2_1
X_18013_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ VPWR VGND _10876_ sg13g2_buf_1
X_18014_ _10876_ _08891_ VPWR VGND _10877_ sg13g2_nand2b_1
X_18015_ _08518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ VPWR VGND _10878_ sg13g2_nor2b_1
X_18016_ _09071_ _10876_ VPWR VGND _10879_ sg13g2_nor2b_1
X_18017_ _08491_ _10874_ _10877_ _10878_ _10879_ VPWR 
+ VGND
+ _10880_ sg13g2_a221oi_1
X_18018_ _10873_ _10875_ _10880_ VPWR VGND _10881_ sg13g2_nor3_1
X_18019_ _10875_ _10880_ _10873_ VPWR VGND _10882_ sg13g2_o21ai_1
X_18020_ _08487_ _10881_ _10882_ VPWR VGND _10883_ sg13g2_o21ai_1
X_18021_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[43]\ VPWR VGND _10884_ sg13g2_buf_1
X_18022_ _10809_ VPWR VGND _10885_ sg13g2_buf_1
X_18023_ _08514_ _10885_ VPWR VGND _10886_ sg13g2_and2_1
X_18024_ _08469_ _10810_ VPWR VGND _10887_ sg13g2_xnor2_1
X_18025_ _08468_ _10887_ _08907_ VPWR VGND _10888_ sg13g2_o21ai_1
X_18026_ _08532_ _10887_ VPWR VGND _10889_ sg13g2_nand2_1
X_18027_ _08906_ _10885_ _10889_ VPWR VGND _10890_ sg13g2_o21ai_1
X_18028_ _10885_ _10889_ VPWR VGND _10891_ sg13g2_nor2_1
X_18029_ _10886_ _10888_ _10890_ _08515_ _10891_ VPWR 
+ VGND
+ _10892_ sg13g2_a221oi_1
X_18030_ _10892_ VPWR VGND _10893_ sg13g2_buf_1
X_18031_ _10884_ _10893_ VPWR VGND _10894_ sg13g2_nand2_1
X_18032_ _09061_ _10893_ VPWR VGND _10895_ sg13g2_nand2_1
X_18033_ _08884_ _10871_ VPWR VGND _10896_ sg13g2_nor2_1
X_18034_ _10872_ _10883_ _10894_ _10895_ _10896_ VPWR 
+ VGND
+ _10897_ sg13g2_a221oi_1
X_18035_ _08474_ _10885_ VPWR VGND _10898_ sg13g2_nand2_1
X_18036_ _10885_ _10192_ _10898_ VPWR VGND _10899_ sg13g2_o21ai_1
X_18037_ _08533_ _10887_ VPWR VGND _10900_ sg13g2_nor2_1
X_18038_ _10889_ _10899_ _10900_ VPWR VGND _10901_ sg13g2_a21o_1
X_18039_ _10885_ _10889_ _08508_ VPWR VGND _10902_ sg13g2_nand3b_1
X_18040_ _08578_ _10810_ VPWR VGND _10903_ sg13g2_xor2_1
X_18041_ _09270_ _10903_ _08532_ VPWR VGND _10904_ sg13g2_a21oi_1
X_18042_ _10192_ _10903_ VPWR VGND _10905_ sg13g2_nor2_1
X_18043_ _10904_ _10905_ _10885_ VPWR VGND _10906_ sg13g2_o21ai_1
X_18044_ _08542_ _10902_ _10906_ VPWR VGND _10907_ sg13g2_nand3_1
X_18045_ _08543_ _10901_ _10907_ VPWR VGND _10908_ sg13g2_o21ai_1
X_18046_ _10885_ _10900_ VPWR VGND _10909_ sg13g2_nand2b_1
X_18047_ _08867_ _10811_ _10812_ VPWR VGND _10910_ sg13g2_a21oi_1
X_18048_ _08550_ _10807_ VPWR VGND _10911_ sg13g2_xnor2_1
X_18049_ _10910_ _10911_ VPWR VGND _10912_ sg13g2_xnor2_1
X_18050_ _08549_ _10912_ VPWR VGND _10913_ sg13g2_xnor2_1
X_18051_ _09061_ _10884_ _10893_ VPWR VGND _10914_ sg13g2_nand3_1
X_18052_ _10908_ _10909_ _10913_ _10914_ VPWR VGND 
+ _10915_
+ sg13g2_nand4_1
X_18053_ _10861_ _10862_ VPWR VGND _10916_ sg13g2_xnor2_1
X_18054_ _08605_ _10912_ _10916_ _08921_ VPWR VGND 
+ _10917_
+ sg13g2_a22oi_1
X_18055_ _10897_ _10915_ _10917_ VPWR VGND _10918_ sg13g2_o21ai_1
X_18056_ _08595_ _10802_ VPWR VGND _10919_ sg13g2_and2_1
X_18057_ _10919_ _10803_ VPWR VGND _10920_ sg13g2_nor2_1
X_18058_ _10819_ _10920_ VPWR VGND _10921_ sg13g2_xnor2_1
X_18059_ _08860_ _10921_ VPWR VGND _10922_ sg13g2_nor2_1
X_18060_ _08635_ _10860_ _10870_ _10918_ _10922_ VPWR 
+ VGND
+ _10923_ sg13g2_a221oi_1
X_18061_ _10853_ _10856_ _10858_ _10859_ _10923_ VPWR 
+ VGND
+ _10924_ sg13g2_a221oi_1
X_18062_ _08646_ _10852_ _10924_ VPWR VGND _10925_ sg13g2_nor3_1
X_18063_ _10852_ _10924_ _08646_ VPWR VGND _10926_ sg13g2_o21ai_1
X_18064_ _10844_ _10925_ _10926_ VPWR VGND _10927_ sg13g2_o21ai_1
X_18065_ _10833_ _10842_ VPWR VGND _10928_ sg13g2_nor2_1
X_18066_ _10833_ _10842_ VPWR VGND _10929_ sg13g2_nand2_1
X_18067_ _08843_ _10928_ _10929_ VPWR VGND _10930_ sg13g2_o21ai_1
X_18068_ _10828_ _10930_ VPWR VGND _10931_ sg13g2_xor2_1
X_18069_ _08841_ _10931_ VPWR VGND _10932_ sg13g2_xnor2_1
X_18070_ _08686_ _10931_ VPWR VGND _10933_ sg13g2_xnor2_1
X_18071_ _08940_ _10798_ VPWR VGND _10934_ sg13g2_xor2_1
X_18072_ _10836_ _10934_ VPWR VGND _10935_ sg13g2_xnor2_1
X_18073_ _10927_ _10932_ _10933_ _08943_ _10935_ VPWR 
+ VGND
+ _10936_ sg13g2_a221oi_1
X_18074_ _10927_ _10932_ _10933_ _08943_ _08955_ VPWR 
+ VGND
+ _10937_ sg13g2_a221oi_1
X_18075_ _08955_ _10935_ VPWR VGND _10938_ sg13g2_nor2_1
X_18076_ _10841_ _10936_ _10937_ _10938_ VPWR VGND 
+ _10939_
+ sg13g2_nor4_1
X_18077_ _08724_ _10797_ VPWR VGND _10940_ sg13g2_nand2_1
X_18078_ _10837_ _10838_ _10940_ VPWR VGND _10941_ sg13g2_o21ai_1
X_18079_ _08725_ _10797_ _10941_ VPWR VGND _10942_ sg13g2_o21ai_1
X_18080_ _10942_ VPWR VGND _10943_ sg13g2_buf_1
X_18081_ _08738_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[17]\ VPWR VGND _10944_ sg13g2_xnor2_1
X_18082_ _10943_ _10944_ VPWR VGND _10945_ sg13g2_xnor2_1
X_18083_ _08716_ _10840_ VPWR VGND _10946_ sg13g2_xnor2_1
X_18084_ _08709_ _10945_ _10946_ _08729_ VPWR VGND 
+ _10947_
+ sg13g2_a22oi_1
X_18085_ _10939_ _10947_ VPWR VGND _10948_ sg13g2_nand2b_1
X_18086_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2643_o\ VPWR VGND _10949_ sg13g2_buf_1
X_18087_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[17]\ VPWR VGND _10950_ sg13g2_inv_1
X_18088_ _10950_ _10943_ _08712_ VPWR VGND _10951_ sg13g2_a21oi_1
X_18089_ _10949_ _10951_ VPWR VGND _10952_ sg13g2_nor2b_1
X_18090_ _10950_ _10949_ _10943_ VPWR VGND _10953_ sg13g2_nor3_1
X_18091_ _10445_ _10945_ VPWR VGND _10954_ sg13g2_nand2_1
X_18092_ _08744_ _10945_ _10954_ VPWR VGND _10955_ sg13g2_o21ai_1
X_18093_ _08759_ _10952_ _10953_ _10955_ VPWR VGND 
+ _10956_
+ sg13g2_nor4_1
X_18094_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2641_o[0]\ VPWR VGND _10957_ sg13g2_buf_1
X_18095_ _10957_ _09151_ VPWR VGND _10958_ sg13g2_nand2_1
X_18096_ _10624_ _08760_ VPWR VGND _10959_ sg13g2_nand2_1
X_18097_ _10948_ _10956_ _10958_ _10959_ VPWR VGND 
+ _00517_
+ sg13g2_a22oi_1
X_18098_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2641_o[1]\ VPWR VGND _10960_ sg13g2_buf_1
X_18099_ _10960_ _09151_ VPWR VGND _10961_ sg13g2_nand2_1
X_18100_ _10794_ _08760_ VPWR VGND _10962_ sg13g2_nand2_1
X_18101_ _10948_ _10956_ _10961_ _10962_ VPWR VGND 
+ _00518_
+ sg13g2_a22oi_1
X_18102_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[16]\ VPWR VGND _10963_ sg13g2_buf_1
X_18103_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[15]\ VPWR VGND _10964_ sg13g2_buf_1
X_18104_ _09205_ _10963_ _10964_ VPWR VGND _10965_ sg13g2_a21oi_1
X_18105_ _09205_ _10963_ _08669_ VPWR VGND _10966_ sg13g2_a21oi_1
X_18106_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[14]\ VPWR VGND _10967_ sg13g2_buf_1
X_18107_ _08653_ _10967_ VPWR VGND _10968_ sg13g2_nand2_1
X_18108_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[13]\ VPWR VGND _10969_ sg13g2_buf_1
X_18109_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[9]\ VPWR VGND _10970_ sg13g2_buf_1
X_18110_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[8]\ VPWR VGND _10971_ sg13g2_buf_1
X_18111_ _08417_ _10971_ VPWR VGND _10972_ sg13g2_nor2_1
X_18112_ _10972_ VPWR VGND _10973_ sg13g2_inv_1
X_18113_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[6]\ VPWR VGND _10974_ sg13g2_buf_1
X_18114_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[7]\ VPWR VGND _10975_ sg13g2_buf_1
X_18115_ _08425_ _10974_ _10975_ VPWR VGND _10976_ sg13g2_a21o_1
X_18116_ _10976_ VPWR VGND _10977_ sg13g2_buf_1
X_18117_ _08425_ _10975_ _10974_ VPWR VGND _10978_ sg13g2_and3_1
X_18118_ _10978_ VPWR VGND _10979_ sg13g2_buf_1
X_18119_ _08469_ _10977_ _10979_ VPWR VGND _10980_ sg13g2_a21o_1
X_18120_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[10]\ VPWR VGND _10981_ sg13g2_buf_1
X_18121_ _08434_ _10981_ _10971_ _08436_ VPWR VGND 
+ _10982_
+ sg13g2_a22oi_1
X_18122_ _10982_ VPWR VGND _10983_ sg13g2_inv_1
X_18123_ _08413_ _10970_ _10973_ _10980_ _10983_ VPWR 
+ VGND
+ _10984_ sg13g2_a221oi_1
X_18124_ _10984_ VPWR VGND _10985_ sg13g2_buf_1
X_18125_ _10970_ VPWR VGND _10986_ sg13g2_inv_1
X_18126_ _08434_ _10981_ VPWR VGND _10987_ sg13g2_nand2_1
X_18127_ _08443_ _10986_ _10987_ VPWR VGND _10988_ sg13g2_nand3_1
X_18128_ _08441_ _10981_ _10988_ VPWR VGND _10989_ sg13g2_o21ai_1
X_18129_ _10989_ VPWR VGND _10990_ sg13g2_buf_1
X_18130_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[12]\ VPWR VGND _10991_ sg13g2_buf_1
X_18131_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[11]\ VPWR VGND _10992_ sg13g2_buf_1
X_18132_ _08454_ _10991_ _10992_ VPWR VGND _10993_ sg13g2_a21oi_1
X_18133_ _10985_ _10990_ _10993_ VPWR VGND _10994_ sg13g2_o21ai_1
X_18134_ _08454_ _10991_ _08407_ VPWR VGND _10995_ sg13g2_a21oi_1
X_18135_ _10985_ _10990_ _10995_ VPWR VGND _10996_ sg13g2_o21ai_1
X_18136_ _08454_ _10991_ VPWR VGND _10997_ sg13g2_nand2_1
X_18137_ _08406_ _10992_ VPWR VGND _10998_ sg13g2_nor2_1
X_18138_ _08454_ _10991_ VPWR VGND _10999_ sg13g2_nor2_1
X_18139_ _10997_ _10998_ _10999_ VPWR VGND _11000_ sg13g2_a21oi_1
X_18140_ _10994_ _10996_ _11000_ VPWR VGND _11001_ sg13g2_and3_1
X_18141_ _11001_ VPWR VGND _11002_ sg13g2_buf_1
X_18142_ _10969_ _11002_ VPWR VGND _11003_ sg13g2_nand2_1
X_18143_ _10969_ _11002_ _08463_ VPWR VGND _11004_ sg13g2_o21ai_1
X_18144_ _10968_ _11003_ _11004_ VPWR VGND _11005_ sg13g2_nand3_1
X_18145_ _08653_ _10967_ _11005_ VPWR VGND _11006_ sg13g2_o21ai_1
X_18146_ _11006_ VPWR VGND _11007_ sg13g2_buf_1
X_18147_ _10965_ _10966_ _11007_ VPWR VGND _11008_ sg13g2_o21ai_1
X_18148_ _08725_ _10963_ VPWR VGND _11009_ sg13g2_nand2_1
X_18149_ _08669_ _10964_ VPWR VGND _11010_ sg13g2_nor2_1
X_18150_ _08725_ _10963_ VPWR VGND _11011_ sg13g2_nor2_1
X_18151_ _11009_ _11010_ _11011_ VPWR VGND _11012_ sg13g2_a21oi_1
X_18152_ _11008_ _11012_ VPWR VGND _11013_ sg13g2_nand2_1
X_18153_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2646_o\ VPWR VGND _11014_ sg13g2_buf_1
X_18154_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[17]\ VPWR VGND _11015_ sg13g2_buf_1
X_18155_ _11014_ _08758_ _11015_ VPWR VGND _11016_ sg13g2_o21ai_1
X_18156_ _11015_ _11013_ VPWR VGND _11017_ sg13g2_nand2b_1
X_18157_ _11013_ _11016_ _11017_ VPWR VGND _11018_ sg13g2_o21ai_1
X_18158_ _08712_ _11014_ _08758_ VPWR VGND _11019_ sg13g2_nor3_1
X_18159_ _11015_ _11013_ VPWR VGND _11020_ sg13g2_xor2_1
X_18160_ _08750_ _11019_ _11020_ VPWR VGND _11021_ sg13g2_nor3_1
X_18161_ _08750_ _11018_ _11021_ VPWR VGND _11022_ sg13g2_a21oi_1
X_18162_ _08940_ _10964_ VPWR VGND _11023_ sg13g2_xor2_1
X_18163_ _11007_ _11023_ VPWR VGND _11024_ sg13g2_xnor2_1
X_18164_ _08680_ _11024_ VPWR VGND _11025_ sg13g2_and2_1
X_18165_ _11003_ _11004_ VPWR VGND _11026_ sg13g2_nand2_1
X_18166_ _08682_ _10967_ VPWR VGND _11027_ sg13g2_xor2_1
X_18167_ _11026_ _11027_ VPWR VGND _11028_ sg13g2_xnor2_1
X_18168_ _08463_ _10969_ VPWR VGND _11029_ sg13g2_xnor2_1
X_18169_ _11002_ _11029_ VPWR VGND _11030_ sg13g2_xnor2_1
X_18170_ _10985_ _10990_ VPWR VGND _11031_ sg13g2_nor2_1
X_18171_ _10992_ _11031_ _08617_ VPWR VGND _11032_ sg13g2_a21oi_1
X_18172_ _10992_ _11031_ VPWR VGND _11033_ sg13g2_nor2_1
X_18173_ _11032_ _11033_ VPWR VGND _11034_ sg13g2_nor2_1
X_18174_ _10991_ _08612_ VPWR VGND _11035_ sg13g2_xor2_1
X_18175_ _11034_ _11035_ VPWR VGND _11036_ sg13g2_xnor2_1
X_18176_ _11030_ _11036_ VPWR VGND _11037_ sg13g2_nand2b_1
X_18177_ _08646_ _11036_ VPWR VGND _11038_ sg13g2_nand2_1
X_18178_ _08616_ _10992_ VPWR VGND _11039_ sg13g2_xnor2_1
X_18179_ _11031_ _11039_ VPWR VGND _11040_ sg13g2_xnor2_1
X_18180_ _08578_ _08468_ VPWR VGND _11041_ sg13g2_xor2_1
X_18181_ _08514_ _10974_ VPWR VGND _11042_ sg13g2_and2_1
X_18182_ _10975_ _11042_ VPWR VGND _11043_ sg13g2_xnor2_1
X_18183_ _11041_ _11043_ VPWR VGND _11044_ sg13g2_xnor2_1
X_18184_ _08551_ _10971_ VPWR VGND _11045_ sg13g2_xor2_1
X_18185_ _10980_ _11045_ VPWR VGND _11046_ sg13g2_xnor2_1
X_18186_ _08549_ _11046_ VPWR VGND _11047_ sg13g2_xnor2_1
X_18187_ _08884_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ VPWR VGND _11048_ sg13g2_nand2_1
X_18188_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[60]\ VPWR VGND _11049_ sg13g2_inv_1
X_18189_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[59]\ VPWR VGND _11050_ sg13g2_buf_1
X_18190_ _08889_ _11050_ VPWR VGND _11051_ sg13g2_nor2_1
X_18191_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[58]\ VPWR VGND _11052_ sg13g2_buf_1
X_18192_ _11052_ _09071_ VPWR VGND _11053_ sg13g2_nand2b_1
X_18193_ _08894_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ VPWR VGND _11054_ sg13g2_nor2b_1
X_18194_ _09071_ _11052_ VPWR VGND _11055_ sg13g2_nor2b_1
X_18195_ _08889_ _11050_ _11053_ _11054_ _11055_ VPWR 
+ VGND
+ _11056_ sg13g2_a221oi_1
X_18196_ _11049_ _11051_ _11056_ VPWR VGND _11057_ sg13g2_nor3_1
X_18197_ _11051_ _11056_ _11049_ VPWR VGND _11058_ sg13g2_o21ai_1
X_18198_ _08487_ _11057_ _11058_ VPWR VGND _11059_ sg13g2_o21ai_1
X_18199_ _10975_ _11041_ VPWR VGND _11060_ sg13g2_xnor2_1
X_18200_ _08542_ _10974_ VPWR VGND _11061_ sg13g2_nor2_1
X_18201_ _11042_ _11060_ _11061_ VPWR VGND _11062_ sg13g2_a21oi_1
X_18202_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[62]\ VPWR VGND _11063_ sg13g2_inv_1
X_18203_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ VPWR VGND _11064_ sg13g2_inv_1
X_18204_ _08878_ _11063_ _11064_ _08883_ VPWR VGND 
+ _11065_
+ sg13g2_a22oi_1
X_18205_ _08907_ _11062_ _11065_ VPWR VGND _11066_ sg13g2_o21ai_1
X_18206_ _11048_ _11059_ _11066_ VPWR VGND _11067_ sg13g2_a21o_1
X_18207_ _10974_ _08901_ VPWR VGND _11068_ sg13g2_xnor2_1
X_18208_ _08879_ _11063_ _11068_ VPWR VGND _11069_ sg13g2_o21ai_1
X_18209_ _08907_ _11062_ _11069_ VPWR VGND _11070_ sg13g2_o21ai_1
X_18210_ _11044_ _11047_ _11067_ _11070_ VPWR VGND 
+ _11071_
+ sg13g2_nand4_1
X_18211_ _08868_ _10979_ VPWR VGND _11072_ sg13g2_nor2_1
X_18212_ _08868_ _11043_ _11072_ VPWR VGND _11073_ sg13g2_a21oi_1
X_18213_ _10971_ _09792_ VPWR VGND _11074_ sg13g2_xnor2_1
X_18214_ _08868_ _10977_ _11074_ VPWR VGND _11075_ sg13g2_nor3_1
X_18215_ _11073_ _11074_ _11075_ VPWR VGND _11076_ sg13g2_a21o_1
X_18216_ _08584_ _10970_ VPWR VGND _11077_ sg13g2_xnor2_1
X_18217_ _08550_ _10971_ _10977_ _08578_ _10979_ VPWR 
+ VGND
+ _11078_ sg13g2_a221oi_1
X_18218_ _11078_ VPWR VGND _11079_ sg13g2_buf_1
X_18219_ _10972_ _11079_ VPWR VGND _11080_ sg13g2_nor2_1
X_18220_ _11077_ _11080_ VPWR VGND _11081_ sg13g2_nand2b_1
X_18221_ _10972_ _11079_ _11077_ VPWR VGND _11082_ sg13g2_o21ai_1
X_18222_ _11081_ _11082_ _08577_ VPWR VGND _11083_ sg13g2_a21oi_1
X_18223_ _08605_ _11046_ _11076_ _08534_ _11083_ VPWR 
+ VGND
+ _11084_ sg13g2_a221oi_1
X_18224_ _08861_ _10970_ VPWR VGND _11085_ sg13g2_nand2_1
X_18225_ _08577_ _11080_ _11085_ VPWR VGND _11086_ sg13g2_a21oi_1
X_18226_ _10981_ _08623_ VPWR VGND _11087_ sg13g2_xor2_1
X_18227_ _11081_ _11087_ VPWR VGND _11088_ sg13g2_nand2_1
X_18228_ _10972_ _11079_ _10986_ VPWR VGND _11089_ sg13g2_o21ai_1
X_18229_ _08861_ _08626_ _11089_ VPWR VGND _11090_ sg13g2_a21o_1
X_18230_ _10986_ _10972_ _11079_ VPWR VGND _11091_ sg13g2_nor3_1
X_18231_ _11091_ _10044_ VPWR VGND _11092_ sg13g2_nand2b_1
X_18232_ _11087_ _11090_ _11092_ VPWR VGND _11093_ sg13g2_nand3b_1
X_18233_ _11086_ _11088_ _11093_ VPWR VGND _11094_ sg13g2_o21ai_1
X_18234_ _08615_ _11040_ _11071_ _11084_ _11094_ VPWR 
+ VGND
+ _11095_ sg13g2_a221oi_1
X_18235_ _08861_ _11091_ _11089_ VPWR VGND _11096_ sg13g2_o21ai_1
X_18236_ _08595_ _10981_ VPWR VGND _11097_ sg13g2_xnor2_1
X_18237_ _11096_ _11097_ VPWR VGND _11098_ sg13g2_xnor2_1
X_18238_ _09048_ _11098_ VPWR VGND _11099_ sg13g2_nand2_1
X_18239_ _08615_ _11040_ _11099_ VPWR VGND _11100_ sg13g2_a21oi_1
X_18240_ _08930_ _11040_ VPWR VGND _11101_ sg13g2_nor2_1
X_18241_ _11095_ _11100_ _11101_ VPWR VGND _11102_ sg13g2_nor3_1
X_18242_ _11037_ _11038_ _11102_ VPWR VGND _11103_ sg13g2_a21oi_1
X_18243_ _10999_ _10997_ VPWR VGND _11104_ sg13g2_nor2b_1
X_18244_ _11034_ _11104_ VPWR VGND _11105_ sg13g2_xnor2_1
X_18245_ _08854_ _11105_ VPWR VGND _11106_ sg13g2_nand2_1
X_18246_ _08844_ _11030_ _11106_ VPWR VGND _11107_ sg13g2_a21oi_1
X_18247_ _08844_ _11030_ VPWR VGND _11108_ sg13g2_nor2_1
X_18248_ _11103_ _11107_ _11108_ VPWR VGND _11109_ sg13g2_or3_1
X_18249_ _09720_ _11028_ VPWR VGND _11110_ sg13g2_xnor2_1
X_18250_ _08943_ _11028_ _11109_ _11110_ VPWR VGND 
+ _11111_
+ sg13g2_a22oi_1
X_18251_ _11024_ _08955_ VPWR VGND _11112_ sg13g2_nand2b_1
X_18252_ _11025_ _11111_ _11112_ VPWR VGND _11113_ sg13g2_o21ai_1
X_18253_ _10964_ VPWR VGND _11114_ sg13g2_inv_1
X_18254_ _11114_ _11007_ _08696_ VPWR VGND _11115_ sg13g2_o21ai_1
X_18255_ _11114_ _11007_ VPWR VGND _11116_ sg13g2_nand2_1
X_18256_ _11115_ _11116_ VPWR VGND _11117_ sg13g2_nand2_1
X_18257_ _10963_ _11117_ VPWR VGND _11118_ sg13g2_xor2_1
X_18258_ _08704_ _11118_ VPWR VGND _11119_ sg13g2_xor2_1
X_18259_ _08716_ _11118_ VPWR VGND _11120_ sg13g2_xnor2_1
X_18260_ _11113_ _11119_ _11120_ _08729_ VPWR VGND 
+ _11121_
+ sg13g2_a22oi_1
X_18261_ _11022_ _11121_ VPWR VGND _11122_ sg13g2_nor2_1
X_18262_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2644_o[0]\ VPWR VGND _11123_ sg13g2_buf_1
X_18263_ _08822_ _11014_ VPWR VGND _11124_ sg13g2_nand2_1
X_18264_ _08712_ _11015_ _11014_ VPWR VGND _11125_ sg13g2_nand3_1
X_18265_ _08739_ _11015_ VPWR VGND _11126_ sg13g2_or2_1
X_18266_ _11125_ _11126_ _11013_ VPWR VGND _11127_ sg13g2_mux2_1
X_18267_ _11020_ _11124_ _11127_ VPWR VGND _11128_ sg13g2_o21ai_1
X_18268_ _08709_ _11128_ VPWR VGND _11129_ sg13g2_nand2_1
X_18269_ _11123_ _08977_ _11129_ VPWR VGND _11130_ sg13g2_nand3_1
X_18270_ _10957_ _10619_ VPWR VGND _11131_ sg13g2_nand2_1
X_18271_ _11122_ _11130_ _11131_ VPWR VGND _00519_ sg13g2_o21ai_1
X_18272_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2644_o[1]\ VPWR VGND _11132_ sg13g2_buf_1
X_18273_ _11132_ _08977_ _11129_ VPWR VGND _11133_ sg13g2_nand3_1
X_18274_ _10960_ _10619_ VPWR VGND _11134_ sg13g2_nand2_1
X_18275_ _11122_ _11133_ _11134_ VPWR VGND _00520_ sg13g2_o21ai_1
X_18276_ _08756_ VPWR VGND _11135_ sg13g2_inv_1
X_18277_ _11123_ _10628_ VPWR VGND _11136_ sg13g2_nand2_1
X_18278_ _11135_ _08981_ _11136_ VPWR VGND _11137_ sg13g2_o21ai_1
X_18279_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[16]\ VPWR VGND _11138_ sg13g2_buf_1
X_18280_ _08724_ _11138_ VPWR VGND _11139_ sg13g2_or2_1
X_18281_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[13]\ VPWR VGND _11140_ sg13g2_buf_1
X_18282_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[12]\ VPWR VGND _11141_ sg13g2_buf_1
X_18283_ _08609_ _11141_ VPWR VGND _11142_ sg13g2_nand2_1
X_18284_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[14]\ VPWR VGND _11143_ sg13g2_buf_1
X_18285_ _08650_ _11143_ VPWR VGND _11144_ sg13g2_nand2_1
X_18286_ _11142_ _11144_ VPWR VGND _11145_ sg13g2_nand2_1
X_18287_ _11140_ _11145_ VPWR VGND _11146_ sg13g2_nor2_1
X_18288_ _08462_ _11145_ VPWR VGND _11147_ sg13g2_nor2_1
X_18289_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[9]\ VPWR VGND _11148_ sg13g2_buf_1
X_18290_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[8]\ VPWR VGND _11149_ sg13g2_buf_1
X_18291_ _08416_ _11149_ VPWR VGND _11150_ sg13g2_nor2_1
X_18292_ _11150_ VPWR VGND _11151_ sg13g2_inv_1
X_18293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[6]\ VPWR VGND _11152_ sg13g2_buf_1
X_18294_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[7]\ VPWR VGND _11153_ sg13g2_buf_1
X_18295_ _08425_ _11152_ _11153_ VPWR VGND _11154_ sg13g2_a21o_1
X_18296_ _11154_ VPWR VGND _11155_ sg13g2_buf_1
X_18297_ _08425_ _11153_ _11152_ VPWR VGND _11156_ sg13g2_and3_1
X_18298_ _11156_ VPWR VGND _11157_ sg13g2_buf_1
X_18299_ _08422_ _11155_ _11157_ VPWR VGND _11158_ sg13g2_a21o_1
X_18300_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[10]\ VPWR VGND _11159_ sg13g2_buf_1
X_18301_ _08433_ _11159_ _11149_ _08417_ VPWR VGND 
+ _11160_
+ sg13g2_a22oi_1
X_18302_ _11160_ VPWR VGND _11161_ sg13g2_inv_1
X_18303_ _08412_ _11148_ _11151_ _11158_ _11161_ VPWR 
+ VGND
+ _11162_ sg13g2_a221oi_1
X_18304_ _11162_ VPWR VGND _11163_ sg13g2_buf_1
X_18305_ _08433_ _11159_ VPWR VGND _11164_ sg13g2_nand2_1
X_18306_ _08412_ _11148_ VPWR VGND _11165_ sg13g2_nor2_1
X_18307_ _08433_ _11159_ VPWR VGND _11166_ sg13g2_nor2_1
X_18308_ _11164_ _11165_ _11166_ VPWR VGND _11167_ sg13g2_a21o_1
X_18309_ _11167_ VPWR VGND _11168_ sg13g2_buf_1
X_18310_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[11]\ VPWR VGND _11169_ sg13g2_inv_1
X_18311_ _11163_ _11168_ _11169_ VPWR VGND _11170_ sg13g2_o21ai_1
X_18312_ _11163_ _11168_ _08639_ VPWR VGND _11171_ sg13g2_o21ai_1
X_18313_ _08609_ _11141_ VPWR VGND _11172_ sg13g2_or2_1
X_18314_ _08639_ _11169_ VPWR VGND _11173_ sg13g2_nand2_1
X_18315_ _11170_ _11171_ _11172_ _11173_ VPWR VGND 
+ _11174_
+ sg13g2_nand4_1
X_18316_ _11174_ VPWR VGND _11175_ sg13g2_buf_1
X_18317_ _11146_ _11147_ _11175_ VPWR VGND _11176_ sg13g2_o21ai_1
X_18318_ _08462_ _11140_ VPWR VGND _11177_ sg13g2_nor2_1
X_18319_ _08651_ _11143_ VPWR VGND _11178_ sg13g2_nor2_1
X_18320_ _11144_ _11177_ _11178_ VPWR VGND _11179_ sg13g2_a21oi_1
X_18321_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[15]\ VPWR VGND _11180_ sg13g2_buf_1
X_18322_ _11176_ _11179_ _11180_ VPWR VGND _11181_ sg13g2_a21oi_1
X_18323_ _11180_ _11176_ _11179_ VPWR VGND _11182_ sg13g2_nand3_1
X_18324_ _08696_ _11181_ _11182_ VPWR VGND _11183_ sg13g2_o21ai_1
X_18325_ _08724_ _11138_ VPWR VGND _11184_ sg13g2_and2_1
X_18326_ _11139_ _11183_ _11184_ VPWR VGND _11185_ sg13g2_a21o_1
X_18327_ _11185_ VPWR VGND _11186_ sg13g2_buf_1
X_18328_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[17]\ VPWR VGND _11187_ sg13g2_buf_1
X_18329_ _08738_ _11187_ VPWR VGND _11188_ sg13g2_xor2_1
X_18330_ _11186_ _11188_ VPWR VGND _11189_ sg13g2_xnor2_1
X_18331_ _08708_ _11189_ VPWR VGND _11190_ sg13g2_and2_1
X_18332_ _08741_ _11189_ VPWR VGND _11191_ sg13g2_or2_1
X_18333_ _08742_ _11189_ VPWR VGND _11192_ sg13g2_nand2_1
X_18334_ _08650_ _11143_ VPWR VGND _11193_ sg13g2_xor2_1
X_18335_ _11193_ VPWR VGND _11194_ sg13g2_buf_1
X_18336_ _11140_ _11194_ VPWR VGND _11195_ sg13g2_nand2_1
X_18337_ _08463_ _11194_ VPWR VGND _11196_ sg13g2_nand2_1
X_18338_ _11195_ _11196_ _11175_ VPWR VGND _11197_ sg13g2_a21o_1
X_18339_ _08455_ _11141_ VPWR VGND _11198_ sg13g2_and2_1
X_18340_ _11198_ VPWR VGND _11199_ sg13g2_buf_1
X_18341_ _11140_ _11199_ _11194_ VPWR VGND _11200_ sg13g2_nor3_1
X_18342_ _08660_ _11199_ _11194_ VPWR VGND _11201_ sg13g2_nor3_1
X_18343_ _11200_ _11201_ _11175_ VPWR VGND _11202_ sg13g2_o21ai_1
X_18344_ _11140_ _11199_ _11194_ VPWR VGND _11203_ sg13g2_nand3_1
X_18345_ _08660_ _11199_ _11194_ VPWR VGND _11204_ sg13g2_nand3_1
X_18346_ _08660_ _11140_ _11194_ VPWR VGND _11205_ sg13g2_nand3_1
X_18347_ _08462_ _11140_ _11194_ VPWR VGND _11206_ sg13g2_or3_1
X_18348_ _11203_ _11204_ _11205_ _11206_ VPWR VGND 
+ _11207_
+ sg13g2_and4_1
X_18349_ _11197_ _11202_ _11207_ VPWR VGND _11208_ sg13g2_nand3_1
X_18350_ _11208_ VPWR VGND _11209_ sg13g2_buf_1
X_18351_ _11159_ _08623_ VPWR VGND _11210_ sg13g2_xnor2_1
X_18352_ _11148_ VPWR VGND _11211_ sg13g2_inv_1
X_18353_ _08436_ _11149_ _11155_ _08469_ _11157_ VPWR 
+ VGND
+ _11212_ sg13g2_a221oi_1
X_18354_ _11212_ VPWR VGND _11213_ sg13g2_buf_1
X_18355_ _11211_ _11150_ _11213_ VPWR VGND _11214_ sg13g2_nor3_1
X_18356_ _11150_ _11213_ _11211_ VPWR VGND _11215_ sg13g2_o21ai_1
X_18357_ _08576_ _11214_ _11215_ VPWR VGND _11216_ sg13g2_o21ai_1
X_18358_ _08576_ _11215_ VPWR VGND _11217_ sg13g2_nor2_1
X_18359_ _08625_ _11216_ _11217_ VPWR VGND _11218_ sg13g2_a21oi_1
X_18360_ _08582_ _11148_ VPWR VGND _11219_ sg13g2_xnor2_1
X_18361_ _11150_ _11213_ _11219_ VPWR VGND _11220_ sg13g2_nor3_1
X_18362_ _11150_ _11213_ VPWR VGND _11221_ sg13g2_nor2_1
X_18363_ _08583_ _11148_ VPWR VGND _11222_ sg13g2_nand2_1
X_18364_ _08576_ _11221_ _11222_ VPWR VGND _11223_ sg13g2_a21oi_1
X_18365_ _11210_ _11220_ _11223_ VPWR VGND _11224_ sg13g2_nor3_1
X_18366_ _11210_ _11218_ _11224_ VPWR VGND _11225_ sg13g2_a21o_1
X_18367_ _11221_ _11219_ VPWR VGND _11226_ sg13g2_xnor2_1
X_18368_ _08550_ _11149_ VPWR VGND _11227_ sg13g2_xor2_1
X_18369_ _11158_ _11227_ VPWR VGND _11228_ sg13g2_xnor2_1
X_18370_ _08604_ _11228_ VPWR VGND _11229_ sg13g2_nand2_1
X_18371_ _08576_ _11226_ _11229_ VPWR VGND _11230_ sg13g2_o21ai_1
X_18372_ _11149_ _09792_ VPWR VGND _11231_ sg13g2_xnor2_1
X_18373_ _11157_ _11231_ VPWR VGND _11232_ sg13g2_and2_1
X_18374_ _11155_ _11231_ VPWR VGND _11233_ sg13g2_nor2_1
X_18375_ _11232_ _11233_ _11041_ VPWR VGND _11234_ sg13g2_o21ai_1
X_18376_ _08867_ _08468_ _11231_ VPWR VGND _11235_ sg13g2_and3_1
X_18377_ _08867_ _08468_ _11231_ VPWR VGND _11236_ sg13g2_nor3_1
X_18378_ _08513_ _11152_ VPWR VGND _11237_ sg13g2_nand2_1
X_18379_ _11153_ _11237_ VPWR VGND _11238_ sg13g2_xnor2_1
X_18380_ _11235_ _11236_ _11238_ VPWR VGND _11239_ sg13g2_o21ai_1
X_18381_ _08542_ _11152_ VPWR VGND _11240_ sg13g2_or2_1
X_18382_ _11234_ _11239_ _11240_ _11237_ _08907_ VPWR 
+ VGND
+ _11241_ sg13g2_a221oi_1
X_18383_ _08548_ _11228_ VPWR VGND _11242_ sg13g2_xor2_1
X_18384_ _09361_ _11238_ VPWR VGND _11243_ sg13g2_xnor2_1
X_18385_ _08872_ _11242_ _11243_ VPWR VGND _11244_ sg13g2_nor3_1
X_18386_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ VPWR VGND _11245_ sg13g2_buf_1
X_18387_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ VPWR VGND _11246_ sg13g2_buf_1
X_18388_ _11246_ _08489_ VPWR VGND _11247_ sg13g2_nand2b_1
X_18389_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ VPWR VGND _11248_ sg13g2_buf_1
X_18390_ _11248_ _08498_ VPWR VGND _11249_ sg13g2_nor2b_1
X_18391_ _08494_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ VPWR VGND _11250_ sg13g2_nand2b_1
X_18392_ _08498_ _11248_ VPWR VGND _11251_ sg13g2_nand2b_1
X_18393_ _11249_ _11250_ _11251_ VPWR VGND _11252_ sg13g2_o21ai_1
X_18394_ _08489_ _11246_ VPWR VGND _11253_ sg13g2_nor2b_1
X_18395_ _08486_ _11245_ _11247_ _11252_ _11253_ VPWR 
+ VGND
+ _11254_ sg13g2_a221oi_1
X_18396_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ VPWR VGND _11255_ sg13g2_buf_1
X_18397_ _11255_ _08882_ VPWR VGND _11256_ sg13g2_nand2b_1
X_18398_ _08486_ _11245_ _11256_ VPWR VGND _11257_ sg13g2_o21ai_1
X_18399_ _08482_ _11255_ VPWR VGND _11258_ sg13g2_nand2_1
X_18400_ _11254_ _11257_ _11258_ VPWR VGND _11259_ sg13g2_o21ai_1
X_18401_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[81]\ VPWR VGND _11260_ sg13g2_inv_1
X_18402_ _08878_ _11260_ VPWR VGND _11261_ sg13g2_nand2_1
X_18403_ _11152_ _08901_ VPWR VGND _11262_ sg13g2_xnor2_1
X_18404_ _08878_ _11260_ _11262_ VPWR VGND _11263_ sg13g2_o21ai_1
X_18405_ _11234_ _11239_ _11259_ _11261_ _11263_ VPWR 
+ VGND
+ _11264_ sg13g2_a221oi_1
X_18406_ _11230_ _11241_ _11244_ _11264_ VPWR VGND 
+ _11265_
+ sg13g2_nor4_1
X_18407_ _08584_ _11214_ _11215_ VPWR VGND _11266_ sg13g2_o21ai_1
X_18408_ _11166_ _11164_ VPWR VGND _11267_ sg13g2_nand2b_1
X_18409_ _11266_ _11267_ VPWR VGND _11268_ sg13g2_xnor2_1
X_18410_ _08589_ _11268_ VPWR VGND _11269_ sg13g2_nand2_1
X_18411_ _11225_ _11265_ _11269_ VPWR VGND _11270_ sg13g2_o21ai_1
X_18412_ _11169_ _11163_ _11168_ VPWR VGND _11271_ sg13g2_nor3_1
X_18413_ _08408_ _11271_ _11170_ VPWR VGND _11272_ sg13g2_o21ai_1
X_18414_ _08456_ _11141_ VPWR VGND _11273_ sg13g2_xnor2_1
X_18415_ _11272_ _11273_ VPWR VGND _11274_ sg13g2_xnor2_1
X_18416_ _11163_ _11168_ VPWR VGND _11275_ sg13g2_nor2_1
X_18417_ _08616_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[11]\ VPWR VGND _11276_ sg13g2_xor2_1
X_18418_ _11275_ _11276_ VPWR VGND _11277_ sg13g2_xnor2_1
X_18419_ _08568_ _11274_ _11277_ VPWR VGND _11278_ sg13g2_a21o_1
X_18420_ _09106_ _10767_ _11274_ VPWR VGND _11279_ sg13g2_mux2_1
X_18421_ _11270_ _11278_ _11279_ VPWR VGND _11280_ sg13g2_o21ai_1
X_18422_ _08568_ _11274_ _11270_ _11277_ _08635_ VPWR 
+ VGND
+ _11281_ sg13g2_a221oi_1
X_18423_ _08660_ _11140_ VPWR VGND _11282_ sg13g2_xor2_1
X_18424_ _08644_ _11282_ VPWR VGND _11283_ sg13g2_and2_1
X_18425_ _08645_ _11282_ VPWR VGND _11284_ sg13g2_nor2_1
X_18426_ _11175_ _11142_ VPWR VGND _11285_ sg13g2_nand2_1
X_18427_ _11283_ _11284_ _11285_ VPWR VGND _11286_ sg13g2_mux2_1
X_18428_ _09720_ _11286_ VPWR VGND _11287_ sg13g2_or2_1
X_18429_ _11209_ _11280_ _11281_ _11287_ VPWR VGND 
+ _11288_
+ sg13g2_nor4_1
X_18430_ _11286_ _11209_ _09720_ VPWR VGND _11289_ sg13g2_nand3b_1
X_18431_ _11280_ _11281_ _11289_ VPWR VGND _11290_ sg13g2_nor3_1
X_18432_ _08683_ _11209_ VPWR VGND _11291_ sg13g2_nand2_1
X_18433_ _09720_ VPWR VGND _11292_ sg13g2_inv_1
X_18434_ _11197_ _11202_ _11207_ VPWR VGND _11293_ sg13g2_and3_1
X_18435_ _11285_ _11282_ VPWR VGND _11294_ sg13g2_xnor2_1
X_18436_ _11292_ _08646_ _11293_ _11294_ VPWR VGND 
+ _11295_
+ sg13g2_nand4_1
X_18437_ _09720_ _08646_ _11209_ _11294_ VPWR VGND 
+ _11296_
+ sg13g2_nand4_1
X_18438_ _11291_ _11295_ _11296_ VPWR VGND _11297_ sg13g2_nand3_1
X_18439_ _11288_ _11290_ _11297_ VPWR VGND _11298_ sg13g2_nor3_1
X_18440_ _08724_ _11138_ VPWR VGND _11299_ sg13g2_xor2_1
X_18441_ _11183_ _11299_ VPWR VGND _11300_ sg13g2_xnor2_1
X_18442_ _11176_ _11179_ VPWR VGND _11301_ sg13g2_nand2_1
X_18443_ _08669_ _11180_ VPWR VGND _11302_ sg13g2_xnor2_1
X_18444_ _11301_ _11302_ VPWR VGND _11303_ sg13g2_xnor2_1
X_18445_ _08728_ _11300_ _11303_ VPWR VGND _11304_ sg13g2_a21oi_1
X_18446_ _08702_ _10344_ _11300_ VPWR VGND _11305_ sg13g2_mux2_1
X_18447_ _11298_ _11304_ _11305_ VPWR VGND _11306_ sg13g2_a21oi_1
X_18448_ _08728_ _11300_ _08955_ VPWR VGND _11307_ sg13g2_a21oi_1
X_18449_ _08681_ _11304_ _11307_ _11298_ VPWR VGND 
+ _11308_
+ sg13g2_a22oi_1
X_18450_ _11306_ _11308_ VPWR VGND _11309_ sg13g2_nand2_1
X_18451_ _11191_ _11192_ _11309_ VPWR VGND _11310_ sg13g2_a21oi_1
X_18452_ _11187_ _11186_ _08822_ VPWR VGND _11311_ sg13g2_o21ai_1
X_18453_ _11187_ _11186_ VPWR VGND _11312_ sg13g2_nand2_1
X_18454_ _11311_ _11312_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2649_o\ VPWR VGND _11313_ sg13g2_a21oi_1
X_18455_ _08759_ _11313_ VPWR VGND _11314_ sg13g2_nor2_1
X_18456_ _11190_ _11310_ _11314_ VPWR VGND _11315_ sg13g2_o21ai_1
X_18457_ _11137_ _11315_ VPWR VGND _00521_ sg13g2_and2_1
X_18458_ _11132_ VPWR VGND _11316_ sg13g2_inv_1
X_18459_ _08974_ _10285_ VPWR VGND _11317_ sg13g2_nand2_1
X_18460_ _11316_ _08977_ _11317_ VPWR VGND _11318_ sg13g2_o21ai_1
X_18461_ _11315_ _11318_ VPWR VGND _00522_ sg13g2_and2_1
X_18462_ _08733_ VPWR VGND _11319_ sg13g2_inv_1
X_18463_ _08970_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ sg13g2_buf_1
X_18464_ _07930_ _11319_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ VPWR VGND _00523_ sg13g2_a21oi_1
X_18465_ _09895_ _07930_ _08981_ VPWR VGND _11320_ sg13g2_a21oi_1
X_18466_ _09692_ _09154_ _11320_ VPWR VGND _00524_ sg13g2_a21o_1
X_18467_ _07932_ VPWR VGND _11321_ sg13g2_buf_1
X_18468_ _07929_ VPWR VGND _11322_ sg13g2_inv_1
X_18469_ _07931_ VPWR VGND _11323_ sg13g2_buf_1
X_18470_ _10100_ _11322_ _11323_ VPWR VGND _11324_ sg13g2_o21ai_1
X_18471_ _09895_ _11321_ _11324_ VPWR VGND _00525_ sg13g2_o21ai_1
X_18472_ _10100_ VPWR VGND _11325_ sg13g2_inv_1
X_18473_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2673_o\ _11322_ _11323_ VPWR VGND _11326_ sg13g2_o21ai_1
X_18474_ _11325_ _11321_ _11326_ VPWR VGND _00526_ sg13g2_o21ai_1
X_18475_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2676_o\ VPWR VGND _11327_ sg13g2_inv_1
X_18476_ _11327_ _07930_ _08981_ VPWR VGND _11328_ sg13g2_a21oi_1
X_18477_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2673_o\ _09154_ _11328_ VPWR VGND _00527_ sg13g2_a21o_1
X_18478_ _10599_ _11322_ _11323_ VPWR VGND _11329_ sg13g2_o21ai_1
X_18479_ _11327_ _11321_ _11329_ VPWR VGND _00528_ sg13g2_o21ai_1
X_18480_ _10629_ _11322_ _11323_ VPWR VGND _11330_ sg13g2_o21ai_1
X_18481_ _11319_ _11321_ _11330_ VPWR VGND _00529_ sg13g2_o21ai_1
X_18482_ _10949_ _11322_ _11323_ VPWR VGND _11331_ sg13g2_o21ai_1
X_18483_ _10789_ _11321_ _11331_ VPWR VGND _00530_ sg13g2_o21ai_1
X_18484_ _11014_ VPWR VGND _11332_ sg13g2_inv_1
X_18485_ _11332_ _07930_ _08981_ VPWR VGND _11333_ sg13g2_a21oi_1
X_18486_ _10949_ _09154_ _11333_ VPWR VGND _00531_ sg13g2_a21o_1
X_18487_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2649_o\ _11322_ _11323_ VPWR VGND _11334_ sg13g2_o21ai_1
X_18488_ _11332_ _11321_ _11334_ VPWR VGND _00532_ sg13g2_o21ai_1
X_18489_ _08970_ VPWR VGND _11335_ sg13g2_buf_1
X_18490_ _08833_ _07930_ _08981_ VPWR VGND _11336_ sg13g2_a21oi_1
X_18491_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2649_o\ _11335_ _11336_ VPWR VGND _00533_ sg13g2_a21o_1
X_18492_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2655_o\ _11322_ _11323_ VPWR VGND _11337_ sg13g2_o21ai_1
X_18493_ _08833_ _11321_ _11337_ VPWR VGND _00534_ sg13g2_o21ai_1
X_18494_ _09157_ _07930_ VPWR VGND _11338_ sg13g2_nor2b_1
X_18495_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2655_o\ _10619_ VPWR VGND _11339_ sg13g2_nand2_1
X_18496_ _09154_ _11338_ _11339_ VPWR VGND _00535_ sg13g2_o21ai_1
X_18497_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2661_o\ _07930_ VPWR VGND _11340_ sg13g2_nor2b_1
X_18498_ _09157_ _10619_ VPWR VGND _11341_ sg13g2_nand2_1
X_18499_ _09154_ _11340_ _11341_ VPWR VGND _00536_ sg13g2_o21ai_1
X_18500_ _09692_ _07930_ VPWR VGND _11342_ sg13g2_nor2b_1
X_18501_ _10628_ VPWR VGND _11343_ sg13g2_buf_1
X_18502_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2661_o\ _11343_ VPWR VGND _11344_ sg13g2_nand2_1
X_18503_ _09154_ _11342_ _11344_ VPWR VGND _00537_ sg13g2_o21ai_1
X_18504_ \atbs_core_0.analog_trigger_0.counter_value[0]\ VPWR VGND _11345_ sg13g2_buf_1
X_18505_ _11345_ _07680_ VPWR VGND _00538_ sg13g2_xnor2_1
X_18506_ _11345_ _07658_ VPWR VGND _11346_ sg13g2_nand2_1
X_18507_ \atbs_core_0.analog_trigger_0.counter_value[1]\ _11346_ VPWR VGND _00539_ sg13g2_xnor2_1
X_18508_ \atbs_core_0.analog_trigger_0.counter_value[1]\ _11345_ _07657_ VPWR VGND _11347_ sg13g2_nand3_1
X_18509_ _11347_ VPWR VGND _11348_ sg13g2_buf_1
X_18510_ \atbs_core_0.analog_trigger_0.counter_value[2]\ _11348_ VPWR VGND _00540_ sg13g2_xnor2_1
X_18511_ \atbs_core_0.analog_trigger_0.counter_value[2]\ VPWR VGND _11349_ sg13g2_inv_1
X_18512_ \atbs_core_0.analog_trigger_0.period_adj_i[6]\ \atbs_core_0.analog_trigger_0.counter_value[6]\ VPWR VGND _11350_ sg13g2_xnor2_1
X_18513_ \atbs_core_0.analog_trigger_0.counter_value[3]\ VPWR VGND _11351_ sg13g2_buf_1
X_18514_ \atbs_core_0.analog_trigger_0.period_adj_i[3]\ _11351_ VPWR VGND _11352_ sg13g2_xnor2_1
X_18515_ \atbs_core_0.analog_trigger_0.counter_value[5]\ VPWR VGND _11353_ sg13g2_buf_1
X_18516_ \atbs_core_0.analog_trigger_0.period_adj_i[5]\ _11353_ VPWR VGND _11354_ sg13g2_xnor2_1
X_18517_ \atbs_core_0.analog_trigger_0.counter_value[4]\ VPWR VGND _11355_ sg13g2_buf_1
X_18518_ \atbs_core_0.analog_trigger_0.period_adj_i[4]\ _11355_ VPWR VGND _11356_ sg13g2_xnor2_1
X_18519_ _11350_ _11352_ _11354_ _11356_ VPWR VGND 
+ _11357_
+ sg13g2_nand4_1
X_18520_ _11349_ _11348_ _11357_ VPWR VGND _11358_ sg13g2_nor3_1
X_18521_ _11349_ _11348_ VPWR VGND _11359_ sg13g2_nor2_1
X_18522_ _11351_ _11359_ VPWR VGND _11360_ sg13g2_xnor2_1
X_18523_ _11358_ _11360_ VPWR VGND _00541_ sg13g2_nor2_1
X_18524_ _11351_ _11359_ VPWR VGND _11361_ sg13g2_nand2_1
X_18525_ _11355_ _11361_ VPWR VGND _11362_ sg13g2_xor2_1
X_18526_ _11358_ _11362_ VPWR VGND _00542_ sg13g2_nor2_1
X_18527_ _11351_ _11355_ _11359_ VPWR VGND _11363_ sg13g2_nand3_1
X_18528_ _11353_ _11363_ VPWR VGND _11364_ sg13g2_xor2_1
X_18529_ _11358_ _11364_ VPWR VGND _00543_ sg13g2_nor2_1
X_18530_ _11351_ _11355_ _11353_ _11359_ VPWR VGND 
+ _11365_
+ sg13g2_nand4_1
X_18531_ \atbs_core_0.analog_trigger_0.counter_value[6]\ _11365_ VPWR VGND _11366_ sg13g2_xor2_1
X_18532_ _11358_ _11366_ VPWR VGND _00544_ sg13g2_nor2_1
X_18533_ _07734_ _07735_ VPWR VGND _11367_ sg13g2_and2_1
X_18534_ _11367_ VPWR VGND _11368_ sg13g2_buf_1
X_18535_ _11368_ VPWR VGND _11369_ sg13g2_buf_1
X_18536_ _11369_ _08232_ VPWR VGND _11370_ sg13g2_nor2_1
X_18537_ _11370_ VPWR VGND _11371_ sg13g2_buf_1
X_18538_ _07713_ _08197_ _08201_ VPWR VGND _11372_ sg13g2_nand3_1
X_18539_ _11372_ VPWR VGND _11373_ sg13g2_buf_4
X_18540_ _00085_ _11373_ VPWR VGND _11374_ sg13g2_xor2_1
X_18541_ _00087_ VPWR VGND _11375_ sg13g2_buf_1
X_18542_ _11375_ VPWR VGND _11376_ sg13g2_inv_1
X_18543_ _08165_ _08168_ VPWR VGND _11377_ sg13g2_nor2_1
X_18544_ _07788_ _08053_ _07712_ VPWR VGND _11378_ sg13g2_o21ai_1
X_18545_ _11378_ VPWR VGND _11379_ sg13g2_buf_1
X_18546_ _11369_ _07755_ _07788_ _08022_ VPWR VGND 
+ _11380_
+ sg13g2_nor4_1
X_18547_ \atbs_core_0.debouncer_5.debounced\ \atbs_core_0.n1420_q\ _07653_ VPWR VGND _11381_ sg13g2_mux2_1
X_18548_ _11381_ VPWR VGND _11382_ sg13g2_buf_1
X_18549_ _07712_ _11382_ VPWR VGND _11383_ sg13g2_nor2b_1
X_18550_ _11383_ VPWR VGND _11384_ sg13g2_buf_1
X_18551_ _11384_ VPWR VGND _11385_ sg13g2_buf_1
X_18552_ \atbs_core_0.n1406_q[4]\ VPWR VGND _11386_ sg13g2_buf_1
X_18553_ _08162_ _11380_ _11385_ _11386_ VPWR VGND 
+ _11387_
+ sg13g2_a22oi_1
X_18554_ _11377_ _11379_ _11387_ VPWR VGND _11388_ sg13g2_o21ai_1
X_18555_ _11388_ VPWR VGND _11389_ sg13g2_buf_4
X_18556_ _11369_ _08055_ VPWR VGND _11390_ sg13g2_nor2_1
X_18557_ _08133_ _08137_ _11390_ VPWR VGND _11391_ sg13g2_nand3_1
X_18558_ _11391_ VPWR VGND _11392_ sg13g2_buf_1
X_18559_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ VPWR VGND _11393_ sg13g2_buf_1
X_18560_ _00089_ VPWR VGND _11394_ sg13g2_buf_1
X_18561_ \atbs_core_0.n1406_q[3]\ VPWR VGND _11395_ sg13g2_buf_1
X_18562_ _11395_ _11384_ VPWR VGND _11396_ sg13g2_nand2_1
X_18563_ _11369_ _08145_ _11396_ VPWR VGND _11397_ sg13g2_o21ai_1
X_18564_ _11397_ VPWR VGND _11398_ sg13g2_buf_1
X_18565_ _11393_ _11394_ _11398_ VPWR VGND _11399_ sg13g2_and3_1
X_18566_ _11393_ _11379_ VPWR VGND _11400_ sg13g2_nor2_1
X_18567_ _11393_ _11398_ VPWR VGND _11401_ sg13g2_nor2_1
X_18568_ _11392_ _11399_ _11400_ _08139_ _11401_ VPWR 
+ VGND
+ _11402_ sg13g2_a221oi_1
X_18569_ _11376_ _11389_ _11402_ VPWR VGND _11403_ sg13g2_a21o_1
X_18570_ _11403_ VPWR VGND _11404_ sg13g2_buf_2
X_18571_ \atbs_core_0.dac_control_0.dac_counter_value[4]\ VPWR VGND _11405_ sg13g2_buf_1
X_18572_ _11375_ _11405_ VPWR VGND _11406_ sg13g2_nand2_1
X_18573_ _11405_ _11406_ _11389_ VPWR VGND _11407_ sg13g2_mux2_1
X_18574_ _11407_ VPWR VGND _11408_ sg13g2_buf_4
X_18575_ _11371_ _11374_ _11404_ _11408_ VPWR VGND 
+ _11409_
+ sg13g2_nand4_1
X_18576_ \atbs_core_0.dac_control_0.dac_counter_value[6]\ VPWR VGND _11410_ sg13g2_buf_2
X_18577_ _11410_ _11374_ _11404_ _11408_ VPWR VGND 
+ _11411_
+ sg13g2_nand4_1
X_18578_ _11394_ VPWR VGND _11412_ sg13g2_inv_1
X_18579_ _11398_ _11392_ VPWR VGND _11413_ sg13g2_and2_1
X_18580_ _11413_ VPWR VGND _11414_ sg13g2_buf_1
X_18581_ _07728_ _08051_ _08164_ _07744_ _11379_ VPWR 
+ VGND
+ _11415_ sg13g2_a221oi_1
X_18582_ \atbs_core_0.n1406_q[2]\ VPWR VGND _11416_ sg13g2_buf_1
X_18583_ _11416_ _11382_ _07712_ VPWR VGND _11417_ sg13g2_a21oi_1
X_18584_ _08096_ _11415_ _11380_ _08107_ _11417_ VPWR 
+ VGND
+ _11418_ sg13g2_a221oi_1
X_18585_ _11418_ VPWR VGND _11419_ sg13g2_buf_8
X_18586_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ _11419_ VPWR VGND _11420_ sg13g2_xnor2_1
X_18587_ _00079_ VPWR VGND _11421_ sg13g2_buf_1
X_18588_ _11421_ VPWR VGND _11422_ sg13g2_inv_1
X_18589_ \atbs_core_0.n1406_q[1]\ VPWR VGND _11423_ sg13g2_buf_1
X_18590_ _11423_ _11384_ VPWR VGND _11424_ sg13g2_nand2_1
X_18591_ _08065_ _11424_ VPWR VGND _11425_ sg13g2_and2_1
X_18592_ _11425_ VPWR VGND _11426_ sg13g2_buf_1
X_18593_ _11423_ _11382_ _07713_ VPWR VGND _11427_ sg13g2_a21oi_1
X_18594_ _08092_ _11390_ _11426_ _08064_ _11427_ VPWR 
+ VGND
+ _11428_ sg13g2_a221oi_1
X_18595_ _11428_ VPWR VGND _11429_ sg13g2_buf_4
X_18596_ _08013_ _08015_ _11379_ VPWR VGND _11430_ sg13g2_nor3_2
X_18597_ _07789_ _11426_ _07936_ VPWR VGND _11431_ sg13g2_nand3b_1
X_18598_ _11368_ _08022_ _08108_ VPWR VGND _11432_ sg13g2_nor3_1
X_18599_ _07788_ _11432_ _07753_ VPWR VGND _11433_ sg13g2_nand3b_1
X_18600_ _11433_ VPWR VGND _11434_ sg13g2_buf_1
X_18601_ _07713_ _11431_ _11434_ VPWR VGND _11435_ sg13g2_nand3_1
X_18602_ _08090_ _11430_ _11435_ VPWR VGND _11436_ sg13g2_a21oi_1
X_18603_ \atbs_core_0.dac_control_0.dac_counter_value[0]\ VPWR VGND _11437_ sg13g2_buf_1
X_18604_ _11437_ VPWR VGND _11438_ sg13g2_inv_1
X_18605_ _08092_ _11390_ _11438_ VPWR VGND _11439_ sg13g2_a21oi_1
X_18606_ _11369_ _11382_ VPWR VGND _11440_ sg13g2_nand2_1
X_18607_ _11422_ _11437_ _11440_ _11434_ VPWR VGND 
+ _11441_
+ sg13g2_nand4_1
X_18608_ _08090_ _11430_ _11441_ VPWR VGND _11442_ sg13g2_a21oi_1
X_18609_ _11422_ _11429_ _11436_ _11439_ _11442_ VPWR 
+ VGND
+ _11443_ sg13g2_a221oi_1
X_18610_ _00083_ VPWR VGND _11444_ sg13g2_buf_1
X_18611_ _11444_ _11419_ VPWR VGND _11445_ sg13g2_nand2b_1
X_18612_ _11420_ _11443_ _11445_ VPWR VGND _11446_ sg13g2_o21ai_1
X_18613_ _11446_ VPWR VGND _11447_ sg13g2_buf_4
X_18614_ _11412_ _11414_ _11389_ _11376_ _11447_ VPWR 
+ VGND
+ _11448_ sg13g2_a221oi_1
X_18615_ _11448_ VPWR VGND _11449_ sg13g2_buf_2
X_18616_ _11409_ _11411_ _11449_ VPWR VGND _11450_ sg13g2_a21oi_2
X_18617_ _11410_ VPWR VGND _11451_ sg13g2_inv_1
X_18618_ _08232_ _07807_ VPWR VGND _11452_ sg13g2_nand2b_1
X_18619_ _11452_ VPWR VGND _11453_ sg13g2_buf_1
X_18620_ \atbs_core_0.dac_control_0.dac_counter_value[5]\ VPWR VGND _11454_ sg13g2_buf_1
X_18621_ _11454_ VPWR VGND _11455_ sg13g2_inv_1
X_18622_ _11455_ _11373_ VPWR VGND _11456_ sg13g2_or2_1
X_18623_ _11451_ _11453_ _11456_ VPWR VGND _11457_ sg13g2_a21oi_1
X_18624_ _11410_ _11371_ _11457_ VPWR VGND _11458_ sg13g2_a21o_1
X_18625_ _00093_ VPWR VGND _11459_ sg13g2_buf_1
X_18626_ _11459_ VPWR VGND _11460_ sg13g2_inv_1
X_18627_ _07836_ _11369_ spike_o VPWR VGND _11461_ sg13g2_o21ai_1
X_18628_ _11461_ \atbs_core_0.dac_control_0.sync_chain_0.async_i\ VPWR VGND _11462_ sg13g2_nand2b_1
X_18629_ _11462_ VPWR VGND _11463_ sg13g2_buf_2
X_18630_ _11460_ _00094_ _11463_ VPWR VGND _11464_ sg13g2_nor3_1
X_18631_ _11450_ _11458_ _11464_ VPWR VGND _11465_ sg13g2_o21ai_1
X_18632_ _11409_ _11411_ _11449_ VPWR VGND _11466_ sg13g2_a21o_1
X_18633_ _11466_ VPWR VGND _11467_ sg13g2_buf_2
X_18634_ _11410_ _11371_ _11457_ VPWR VGND _11468_ sg13g2_a21oi_1
X_18635_ _11459_ _00094_ _11463_ VPWR VGND _11469_ sg13g2_nor3_1
X_18636_ _11467_ _11468_ _11469_ VPWR VGND _11470_ sg13g2_nand3_1
X_18637_ _11470_ VPWR VGND _11471_ sg13g2_buf_2
X_18638_ _11465_ _11471_ VPWR VGND _11472_ sg13g2_nand2_1
X_18639_ \atbs_core_0.dac_control_0.n1938_q\ VPWR VGND _11473_ sg13g2_buf_4
X_18640_ _08090_ _11430_ _11432_ _08064_ _11385_ VPWR 
+ VGND
+ _11474_ sg13g2_a221oi_1
X_18641_ _11474_ VPWR VGND _11475_ sg13g2_buf_1
X_18642_ _11475_ _11461_ \atbs_core_0.dac_control_0.sync_chain_0.async_i\ VPWR VGND _11476_ sg13g2_o21ai_1
X_18643_ _11473_ _11476_ VPWR VGND _11477_ sg13g2_and2_1
X_18644_ _11472_ _11477_ _11437_ VPWR VGND _11478_ sg13g2_o21ai_1
X_18645_ _11463_ VPWR VGND _11479_ sg13g2_buf_2
X_18646_ _00037_ VPWR VGND _11480_ sg13g2_buf_1
X_18647_ _11480_ _11475_ VPWR VGND _11481_ sg13g2_xnor2_1
X_18648_ _11389_ VPWR VGND _11482_ sg13g2_inv_1
X_18649_ _11376_ _11482_ VPWR VGND _11483_ sg13g2_nand2_1
X_18650_ _11398_ _11392_ VPWR VGND _11484_ sg13g2_nand2_1
X_18651_ _11484_ VPWR VGND _11485_ sg13g2_buf_2
X_18652_ _11480_ VPWR VGND _11486_ sg13g2_inv_1
X_18653_ _08092_ _11390_ _11486_ VPWR VGND _11487_ sg13g2_a21oi_1
X_18654_ _11369_ _11424_ _11426_ _08064_ _11422_ VPWR 
+ VGND
+ _11488_ sg13g2_a221oi_1
X_18655_ _08092_ _11390_ VPWR VGND _11489_ sg13g2_nand2_1
X_18656_ _11421_ _11480_ _11440_ _11434_ VPWR VGND 
+ _11490_
+ sg13g2_nand4_1
X_18657_ _08090_ _11430_ _11490_ VPWR VGND _11491_ sg13g2_a21oi_1
X_18658_ _11436_ _11487_ _11488_ _11489_ _11491_ VPWR 
+ VGND
+ _11492_ sg13g2_a221oi_1
X_18659_ _11492_ VPWR VGND _11493_ sg13g2_buf_1
X_18660_ _11444_ _11419_ VPWR VGND _11494_ sg13g2_nor2_1
X_18661_ _11485_ _11493_ _11494_ VPWR VGND _11495_ sg13g2_nor3_1
X_18662_ _11444_ _11419_ VPWR VGND _11496_ sg13g2_nand2_1
X_18663_ _11412_ _11485_ _11496_ VPWR VGND _11497_ sg13g2_a21oi_1
X_18664_ _11444_ _11419_ _11394_ VPWR VGND _11498_ sg13g2_o21ai_1
X_18665_ _11394_ _11398_ _11392_ VPWR VGND _11499_ sg13g2_nand3_1
X_18666_ _11493_ _11498_ _11499_ VPWR VGND _11500_ sg13g2_o21ai_1
X_18667_ _11495_ _11497_ _11500_ VPWR VGND _11501_ sg13g2_or3_1
X_18668_ _11501_ VPWR VGND _11502_ sg13g2_buf_1
X_18669_ _11375_ _11389_ VPWR VGND _11503_ sg13g2_nand2_1
X_18670_ _11373_ _11503_ VPWR VGND _11504_ sg13g2_nand2_1
X_18671_ _11454_ _11503_ VPWR VGND _11505_ sg13g2_nand2_1
X_18672_ _11455_ _11373_ VPWR VGND _11506_ sg13g2_xnor2_1
X_18673_ _11376_ _11389_ VPWR VGND _11507_ sg13g2_xnor2_1
X_18674_ _11412_ _11414_ VPWR VGND _11508_ sg13g2_xnor2_1
X_18675_ _11444_ _11419_ VPWR VGND _11509_ sg13g2_xnor2_1
X_18676_ _11421_ _11429_ VPWR VGND _11510_ sg13g2_xnor2_1
X_18677_ _11509_ _11481_ _11510_ VPWR VGND _11511_ sg13g2_nor3_1
X_18678_ _11506_ _11507_ _11508_ _11511_ VPWR VGND 
+ _11512_
+ sg13g2_and4_1
X_18679_ _11483_ _11502_ _11504_ _11505_ _11512_ VPWR 
+ VGND
+ _11513_ sg13g2_a221oi_1
X_18680_ _11454_ _11373_ _11453_ VPWR VGND _11514_ sg13g2_a21oi_1
X_18681_ _11513_ _11514_ VPWR VGND _11515_ sg13g2_nor2b_1
X_18682_ _11495_ _11497_ _11500_ VPWR VGND _11516_ sg13g2_nor3_1
X_18683_ _11454_ _11373_ _11482_ _11376_ _11516_ VPWR 
+ VGND
+ _11517_ sg13g2_a221oi_1
X_18684_ _11454_ _11373_ _11503_ VPWR VGND _11518_ sg13g2_a21o_1
X_18685_ _11454_ _11373_ _11518_ VPWR VGND _11519_ sg13g2_o21ai_1
X_18686_ _11371_ _11512_ _11517_ _11519_ VPWR VGND 
+ _11520_
+ sg13g2_or4_1
X_18687_ _11410_ _11460_ VPWR VGND _11521_ sg13g2_nor2_1
X_18688_ _11459_ _11515_ _11520_ _11521_ VPWR VGND 
+ _11522_
+ sg13g2_a22oi_1
X_18689_ _11522_ VPWR VGND _11523_ sg13g2_buf_1
X_18690_ _11473_ VPWR VGND _11524_ sg13g2_inv_1
X_18691_ _11524_ _07805_ VPWR VGND _11525_ sg13g2_nor2_1
X_18692_ _11479_ _11481_ _11523_ _11525_ VPWR VGND 
+ _11526_
+ sg13g2_nand4_1
X_18693_ _11467_ _11468_ VPWR VGND _11527_ sg13g2_nand2_1
X_18694_ _11460_ _11527_ VPWR VGND _11528_ sg13g2_xnor2_1
X_18695_ _07805_ _11461_ VPWR VGND _11529_ sg13g2_nor2_1
X_18696_ _11529_ VPWR VGND _11530_ sg13g2_buf_1
X_18697_ _11438_ _11475_ _11530_ _11525_ VPWR VGND 
+ _11531_
+ sg13g2_and4_1
X_18698_ _00094_ _11528_ _11531_ VPWR VGND _11532_ sg13g2_o21ai_1
X_18699_ _11478_ _11526_ _11532_ VPWR VGND _00552_ sg13g2_nand3_1
X_18700_ \atbs_core_0.dac_control_0.dac_counter_value[1]\ VPWR VGND _11533_ sg13g2_inv_1
X_18701_ _11473_ _07805_ VPWR VGND _11534_ sg13g2_nand2_1
X_18702_ _11465_ _11471_ _11534_ VPWR VGND _11535_ sg13g2_nand3_1
X_18703_ _11535_ VPWR VGND _11536_ sg13g2_buf_4
X_18704_ _11536_ VPWR VGND _11537_ sg13g2_buf_16
X_18705_ _11524_ \atbs_core_0.dac_control_0.dac_init_value[1]\ _11537_ VPWR VGND _11538_ sg13g2_a21oi_2
X_18706_ _11437_ _11480_ _11479_ VPWR VGND _11539_ sg13g2_mux2_1
X_18707_ _11475_ _11539_ VPWR VGND _11540_ sg13g2_nand2_1
X_18708_ _11510_ _11540_ VPWR VGND _11541_ sg13g2_xnor2_1
X_18709_ _11473_ _11541_ VPWR VGND _11542_ sg13g2_and2_1
X_18710_ _11530_ _11523_ _11542_ VPWR VGND _11543_ sg13g2_o21ai_1
X_18711_ _11533_ _11537_ _11538_ _11543_ VPWR VGND 
+ _00553_
+ sg13g2_a22oi_1
X_18712_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ VPWR VGND _11544_ sg13g2_inv_1
X_18713_ _11420_ _11443_ VPWR VGND _11545_ sg13g2_xor2_1
X_18714_ _11465_ _11471_ _11525_ VPWR VGND _11546_ sg13g2_nand3_1
X_18715_ _11546_ VPWR VGND _11547_ sg13g2_buf_2
X_18716_ _11530_ _11545_ _11547_ VPWR VGND _11548_ sg13g2_a21oi_1
X_18717_ _11509_ _11493_ VPWR VGND _11549_ sg13g2_xnor2_1
X_18718_ _11479_ _11523_ _11549_ VPWR VGND _11550_ sg13g2_nand3_1
X_18719_ _11473_ \atbs_core_0.dac_control_0.dac_init_value[2]\ _11537_ VPWR VGND _11551_ sg13g2_nor3_2
X_18720_ _11544_ _11537_ _11548_ _11550_ _11551_ VPWR 
+ VGND
+ _00554_ sg13g2_a221oi_1
X_18721_ _11393_ VPWR VGND _11552_ sg13g2_inv_1
X_18722_ _11493_ _11494_ _11496_ VPWR VGND _11553_ sg13g2_o21ai_1
X_18723_ _11508_ _11553_ VPWR VGND _11554_ sg13g2_xnor2_1
X_18724_ _11479_ _11523_ _11554_ VPWR VGND _11555_ sg13g2_nand3_1
X_18725_ _11393_ _11414_ VPWR VGND _11556_ sg13g2_xnor2_1
X_18726_ _11447_ _11556_ VPWR VGND _11557_ sg13g2_xnor2_1
X_18727_ _11530_ _11557_ _11547_ VPWR VGND _11558_ sg13g2_a21oi_1
X_18728_ _11473_ \atbs_core_0.dac_control_0.dac_init_value[3]\ _11537_ VPWR VGND _11559_ sg13g2_nor3_2
X_18729_ _11552_ _11537_ _11555_ _11558_ _11559_ VPWR 
+ VGND
+ _00555_ sg13g2_a221oi_1
X_18730_ _11405_ VPWR VGND _11560_ sg13g2_inv_1
X_18731_ _11507_ _11502_ VPWR VGND _11561_ sg13g2_xnor2_1
X_18732_ _11479_ _11523_ _11561_ VPWR VGND _11562_ sg13g2_nand3_1
X_18733_ _11552_ _11447_ _11412_ VPWR VGND _11563_ sg13g2_a21oi_1
X_18734_ _11393_ _11447_ VPWR VGND _11564_ sg13g2_nand2_1
X_18735_ _11563_ _11564_ _11485_ VPWR VGND _11565_ sg13g2_mux2_1
X_18736_ _11560_ _11389_ VPWR VGND _11566_ sg13g2_xnor2_1
X_18737_ _11565_ _11566_ VPWR VGND _11567_ sg13g2_xnor2_1
X_18738_ _11530_ _11567_ _11547_ VPWR VGND _11568_ sg13g2_a21oi_1
X_18739_ _11473_ \atbs_core_0.dac_control_0.dac_init_value[4]\ _11537_ VPWR VGND _11569_ sg13g2_nor3_2
X_18740_ _11560_ _11537_ _11562_ _11568_ _11569_ VPWR 
+ VGND
+ _00556_ sg13g2_a221oi_1
X_18741_ _11483_ _11502_ VPWR VGND _11570_ sg13g2_nand2_1
X_18742_ _11503_ _11570_ VPWR VGND _11571_ sg13g2_nand2_1
X_18743_ _11506_ _11571_ VPWR VGND _11572_ sg13g2_xnor2_1
X_18744_ _11479_ _11523_ _11572_ VPWR VGND _11573_ sg13g2_nand3_1
X_18745_ _11404_ _11408_ VPWR VGND _11574_ sg13g2_nand2_1
X_18746_ _11449_ _11574_ VPWR VGND _11575_ sg13g2_nor2_1
X_18747_ _11374_ _11575_ VPWR VGND _11576_ sg13g2_xnor2_1
X_18748_ _11479_ _11576_ _11473_ VPWR VGND _11577_ sg13g2_o21ai_1
X_18749_ _11536_ _11577_ VPWR VGND _11578_ sg13g2_nor2_1
X_18750_ _11473_ \atbs_core_0.dac_control_0.dac_init_value[5]\ _11536_ VPWR VGND _11579_ sg13g2_nor3_1
X_18751_ _11455_ _11537_ _11573_ _11578_ _11579_ VPWR 
+ VGND
+ _00557_ sg13g2_a221oi_1
X_18752_ _11524_ _11537_ VPWR VGND _11580_ sg13g2_nor2_2
X_18753_ _11374_ _11404_ _11408_ VPWR VGND _11581_ sg13g2_nand3_1
X_18754_ _11449_ _11581_ _11456_ VPWR VGND _11582_ sg13g2_o21ai_1
X_18755_ _11410_ _11371_ VPWR VGND _11583_ sg13g2_xnor2_1
X_18756_ _11582_ _11583_ VPWR VGND _11584_ sg13g2_xnor2_1
X_18757_ _11530_ _11584_ VPWR VGND _11585_ sg13g2_nand2_1
X_18758_ _11410_ _11459_ _11371_ _11530_ VPWR VGND 
+ _11586_
+ sg13g2_nor4_1
X_18759_ _11451_ _11459_ _11453_ _11530_ VPWR VGND 
+ _11587_
+ sg13g2_nor4_1
X_18760_ _11517_ _11519_ VPWR VGND _11588_ sg13g2_or2_1
X_18761_ _11588_ VPWR VGND _11589_ sg13g2_buf_1
X_18762_ _11586_ _11587_ _11589_ VPWR VGND _11590_ sg13g2_o21ai_1
X_18763_ _11410_ _11453_ _11479_ VPWR VGND _11591_ sg13g2_nand3_1
X_18764_ _11451_ _11460_ _11371_ _11479_ VPWR VGND 
+ _11592_
+ sg13g2_nand4_1
X_18765_ _11591_ _11592_ _11589_ VPWR VGND _11593_ sg13g2_a21o_1
X_18766_ _11585_ _11590_ _11593_ VPWR VGND _11594_ sg13g2_nand3_1
X_18767_ _11473_ \atbs_core_0.dac_control_0.dac_init_value[6]\ VPWR VGND _11595_ sg13g2_nor2b_1
X_18768_ _11595_ _11410_ _11536_ VPWR VGND _11596_ sg13g2_mux2_1
X_18769_ _11580_ _11594_ _11596_ VPWR VGND _00558_ sg13g2_a21o_1
X_18770_ _11371_ _11589_ _11451_ VPWR VGND _11597_ sg13g2_o21ai_1
X_18771_ _11460_ _11479_ VPWR VGND _11598_ sg13g2_nand2_1
X_18772_ _11371_ _11589_ _11598_ VPWR VGND _11599_ sg13g2_a21oi_1
X_18773_ _11450_ _11458_ _11530_ VPWR VGND _11600_ sg13g2_o21ai_1
X_18774_ _11460_ _11467_ _11468_ _11530_ VPWR VGND 
+ _11601_
+ sg13g2_nand4_1
X_18775_ _11460_ _11600_ _11601_ VPWR VGND _11602_ sg13g2_o21ai_1
X_18776_ _11597_ _11599_ _11602_ VPWR VGND _11603_ sg13g2_a21oi_1
X_18777_ _11524_ \atbs_core_0.dac_control_0.dac_init_value[7]\ VPWR VGND _11604_ sg13g2_nand2_1
X_18778_ \atbs_core_0.dac_control_0.dac_counter_value[7]\ VPWR VGND _11605_ sg13g2_inv_1
X_18779_ _11604_ _11605_ _11536_ VPWR VGND _11606_ sg13g2_mux2_1
X_18780_ _11547_ _11603_ _11606_ VPWR VGND _00559_ sg13g2_o21ai_1
X_18781_ \atbs_core_0.dac_control_0.n1942_q[1]\ \atbs_core_0.dac_control_0.n1942_q[0]\ VPWR VGND _11607_ sg13g2_nand2_1
X_18782_ _00058_ _11607_ VPWR VGND _11608_ sg13g2_or2_1
X_18783_ _07678_ _11524_ _07805_ VPWR VGND _11609_ sg13g2_a21oi_1
X_18784_ \atbs_core_0.dac_control_0.dac_change_in_progress\ _11608_ _11609_ VPWR VGND _00560_ sg13g2_a21o_1
X_18785_ dac_upper_o[0] VPWR VGND _11610_ sg13g2_inv_1
X_18786_ \atbs_core_0.dac_control_0.sync_chain_0.async_i\ _11453_ _11373_ _11482_ VPWR VGND 
+ _11611_
+ sg13g2_and4_1
X_18787_ _11485_ _11611_ VPWR VGND _11612_ sg13g2_and2_1
X_18788_ _11612_ VPWR VGND _11613_ sg13g2_buf_1
X_18789_ _11419_ _11429_ VPWR VGND _11614_ sg13g2_nor2_1
X_18790_ _11475_ _11614_ VPWR VGND _11615_ sg13g2_and2_1
X_18791_ _11610_ _07805_ _11613_ _11615_ VPWR VGND 
+ _00561_
+ sg13g2_a22oi_1
X_18792_ dac_upper_o[1] VPWR VGND _11616_ sg13g2_inv_1
X_18793_ _11429_ _11475_ VPWR VGND _11617_ sg13g2_xnor2_1
X_18794_ _11419_ _11617_ VPWR VGND _11618_ sg13g2_nor2_1
X_18795_ _11616_ _07805_ _11613_ _11618_ VPWR VGND 
+ _00562_
+ sg13g2_a22oi_1
X_18796_ dac_upper_o[2] VPWR VGND _11619_ sg13g2_inv_1
X_18797_ _11475_ _11419_ VPWR VGND _11620_ sg13g2_nor2b_1
X_18798_ _11429_ _11620_ VPWR VGND _11621_ sg13g2_nand2b_1
X_18799_ _11618_ _11621_ VPWR VGND _11622_ sg13g2_nand2b_1
X_18800_ _11619_ _07805_ _11613_ _11622_ VPWR VGND 
+ _00563_
+ sg13g2_a22oi_1
X_18801_ dac_upper_o[3] VPWR VGND _11623_ sg13g2_inv_1
X_18802_ _11419_ _11429_ VPWR VGND _11624_ sg13g2_xnor2_1
X_18803_ _11485_ _11624_ VPWR VGND _11625_ sg13g2_nand2_1
X_18804_ _11485_ _11614_ _11625_ VPWR VGND _11626_ sg13g2_o21ai_1
X_18805_ _11485_ _11615_ VPWR VGND _11627_ sg13g2_nand2_1
X_18806_ _11475_ _11626_ _11627_ VPWR VGND _11628_ sg13g2_o21ai_1
X_18807_ _11623_ _07805_ _11611_ _11628_ VPWR VGND 
+ _00564_
+ sg13g2_a22oi_1
X_18808_ \atbs_core_0.dac_control_1.dac_counter_value[0]\ VPWR VGND _11629_ sg13g2_buf_1
X_18809_ _11629_ VPWR VGND _11630_ sg13g2_inv_1
X_18810_ _08026_ _08051_ _08164_ _08255_ VPWR VGND 
+ _11631_
+ sg13g2_nor4_2
X_18811_ _11369_ _08013_ _08015_ _08257_ VPWR VGND 
+ _11632_
+ sg13g2_or4_1
X_18812_ _11632_ VPWR VGND _11633_ sg13g2_buf_2
X_18813_ _11631_ _11633_ _11440_ VPWR VGND _11634_ sg13g2_o21ai_1
X_18814_ _11634_ VPWR VGND _11635_ sg13g2_buf_1
X_18815_ _00096_ VPWR VGND _11636_ sg13g2_buf_1
X_18816_ _11636_ VPWR VGND _11637_ sg13g2_inv_1
X_18817_ _07713_ _08097_ _08098_ _08293_ VPWR VGND 
+ _11638_
+ sg13g2_and4_1
X_18818_ _07713_ _08295_ _11417_ VPWR VGND _11639_ sg13g2_a21o_1
X_18819_ _08096_ _11638_ _11639_ VPWR VGND _11640_ sg13g2_a21oi_1
X_18820_ _11640_ VPWR VGND _11641_ sg13g2_buf_8
X_18821_ _11637_ _11641_ VPWR VGND _11642_ sg13g2_nand2_1
X_18822_ _08096_ _11638_ _11639_ VPWR VGND _11643_ sg13g2_a21o_1
X_18823_ _11643_ VPWR VGND _11644_ sg13g2_buf_1
X_18824_ _11636_ _11644_ VPWR VGND _11645_ sg13g2_nand2_1
X_18825_ _11630_ _11635_ VPWR VGND _11646_ sg13g2_nand2_1
X_18826_ _07807_ _08260_ _11385_ VPWR VGND _11647_ sg13g2_a21oi_1
X_18827_ _11629_ _11647_ VPWR VGND _11648_ sg13g2_nand2_1
X_18828_ _07715_ _07807_ VPWR VGND _11649_ sg13g2_nand2_1
X_18829_ _07936_ _11649_ VPWR VGND _11650_ sg13g2_nand2_1
X_18830_ _07709_ _07841_ _11650_ VPWR VGND _11651_ sg13g2_o21ai_1
X_18831_ _11651_ VPWR VGND _11652_ sg13g2_buf_1
X_18832_ _00097_ VPWR VGND _11653_ sg13g2_inv_1
X_18833_ spike_o _08269_ _11385_ _11423_ VPWR VGND 
+ _11654_
+ sg13g2_a22oi_1
X_18834_ _08267_ _11426_ _11427_ VPWR VGND _11655_ sg13g2_a21o_1
X_18835_ _08044_ _11654_ _11655_ VPWR VGND _11656_ sg13g2_a21oi_1
X_18836_ _11653_ _11656_ VPWR VGND _11657_ sg13g2_xnor2_1
X_18837_ _08134_ _08135_ _08318_ _11396_ VPWR VGND 
+ _11658_
+ sg13g2_and4_1
X_18838_ _07713_ _08323_ _11385_ _11395_ VPWR VGND 
+ _11659_
+ sg13g2_a22oi_1
X_18839_ _08133_ _11658_ _11659_ VPWR VGND _11660_ sg13g2_a21oi_1
X_18840_ _11660_ VPWR VGND _11661_ sg13g2_buf_2
X_18841_ _00095_ VPWR VGND _11662_ sg13g2_inv_1
X_18842_ _11661_ _11662_ VPWR VGND _11663_ sg13g2_nand2b_1
X_18843_ _00036_ _11652_ _11657_ _11663_ VPWR VGND 
+ _11664_
+ sg13g2_nand4_1
X_18844_ _11642_ _11645_ _11646_ _11648_ _11664_ VPWR 
+ VGND
+ _11665_ sg13g2_a221oi_1
X_18845_ \atbs_core_0.dac_control_1.dac_counter_value[5]\ VPWR VGND _11666_ sg13g2_buf_1
X_18846_ _08195_ _08319_ _07807_ VPWR VGND _11667_ sg13g2_o21ai_1
X_18847_ _11667_ VPWR VGND _11668_ sg13g2_buf_1
X_18848_ _08361_ _11668_ VPWR VGND _11669_ sg13g2_nor2_1
X_18849_ _11666_ _11669_ VPWR VGND _11670_ sg13g2_xnor2_1
X_18850_ _11369_ _08308_ VPWR VGND _11671_ sg13g2_nor2_1
X_18851_ _08165_ _08168_ _11671_ VPWR VGND _11672_ sg13g2_o21ai_1
X_18852_ _11672_ VPWR VGND _11673_ sg13g2_buf_1
X_18853_ _11386_ _11385_ VPWR VGND _11674_ sg13g2_nand2_1
X_18854_ _07713_ _08162_ _08308_ VPWR VGND _11675_ sg13g2_nand3_1
X_18855_ _11674_ _11675_ VPWR VGND _11676_ sg13g2_and2_1
X_18856_ _11676_ VPWR VGND _11677_ sg13g2_buf_1
X_18857_ _00098_ VPWR VGND _11678_ sg13g2_inv_1
X_18858_ _11673_ _11677_ _11678_ VPWR VGND _11679_ sg13g2_a21oi_1
X_18859_ _11678_ _11673_ _11677_ VPWR VGND _11680_ sg13g2_nand3_1
X_18860_ _11679_ _11680_ VPWR VGND _11681_ sg13g2_nor2b_1
X_18861_ _00095_ _11661_ VPWR VGND _11682_ sg13g2_nand2_1
X_18862_ \atbs_core_0.dac_control_1.dac_counter_value[6]\ VPWR VGND _11683_ sg13g2_buf_1
X_18863_ _07734_ _07735_ _08224_ _08319_ _08378_ VPWR 
+ VGND
+ _11684_ sg13g2_a221oi_1
X_18864_ _11684_ VPWR VGND _11685_ sg13g2_buf_1
X_18865_ _11683_ _11685_ VPWR VGND _11686_ sg13g2_xnor2_1
X_18866_ _11670_ _11681_ _11682_ _11686_ VPWR VGND 
+ _11687_
+ sg13g2_and4_1
X_18867_ _08044_ _11654_ _11655_ VPWR VGND _11688_ sg13g2_a21o_1
X_18868_ _11688_ VPWR VGND _11689_ sg13g2_buf_2
X_18869_ _11629_ _11385_ VPWR VGND _11690_ sg13g2_nor2_1
X_18870_ _11631_ _11633_ _11690_ VPWR VGND _11691_ sg13g2_o21ai_1
X_18871_ _11691_ VPWR VGND _11692_ sg13g2_buf_2
X_18872_ _11689_ _11692_ _11653_ VPWR VGND _11693_ sg13g2_o21ai_1
X_18873_ _11693_ VPWR VGND _11694_ sg13g2_buf_1
X_18874_ _11637_ _11644_ _11689_ _11692_ VPWR VGND 
+ _11695_
+ sg13g2_a22oi_1
X_18875_ _11636_ _11641_ _11694_ _11695_ VPWR VGND 
+ _11696_
+ sg13g2_a22oi_1
X_18876_ _11670_ _11681_ _11682_ _11696_ VPWR VGND 
+ _11697_
+ sg13g2_nand4_1
X_18877_ _11697_ VPWR VGND _11698_ sg13g2_buf_2
X_18878_ _08380_ _07807_ VPWR VGND _11699_ sg13g2_nand2b_1
X_18879_ _11699_ VPWR VGND _11700_ sg13g2_buf_1
X_18880_ _00036_ _11652_ VPWR VGND _11701_ sg13g2_nand2_1
X_18881_ _11666_ _08361_ _11668_ VPWR VGND _11702_ sg13g2_nor3_1
X_18882_ _11663_ _11702_ _11679_ VPWR VGND _11703_ sg13g2_nor3_1
X_18883_ _08361_ _11668_ _11666_ VPWR VGND _11704_ sg13g2_o21ai_1
X_18884_ _11702_ _11680_ _11704_ VPWR VGND _11705_ sg13g2_o21ai_1
X_18885_ _11700_ _11701_ _11703_ _11705_ VPWR VGND 
+ _11706_
+ sg13g2_nor4_1
X_18886_ \atbs_core_0.dac_control_1.n2087_q\ VPWR VGND _11707_ sg13g2_buf_1
X_18887_ _11707_ \atbs_core_0.dac_control_1.sync_chain_0.async_i\ VPWR VGND _11708_ sg13g2_nand2_1
X_18888_ _11665_ _11687_ _11698_ _11706_ _11708_ VPWR 
+ VGND
+ _11709_ sg13g2_a221oi_1
X_18889_ _11703_ _11705_ VPWR VGND _11710_ sg13g2_nor2_1
X_18890_ _11683_ _11701_ VPWR VGND _11711_ sg13g2_nor2_1
X_18891_ _11698_ _11710_ _11711_ VPWR VGND _11712_ sg13g2_nand3_1
X_18892_ _11685_ _11711_ VPWR VGND _11713_ sg13g2_nand2_1
X_18893_ _11709_ _11712_ _11713_ VPWR VGND _11714_ sg13g2_and3_1
X_18894_ _11714_ VPWR VGND _11715_ sg13g2_buf_2
X_18895_ _07807_ _08335_ _11385_ _11395_ VPWR VGND 
+ _11716_
+ sg13g2_a22oi_1
X_18896_ _11716_ VPWR VGND _11717_ sg13g2_buf_1
X_18897_ _00095_ _11717_ VPWR VGND _11718_ sg13g2_nor2_1
X_18898_ \atbs_core_0.dac_control_1.dac_counter_value[2]\ VPWR VGND _11719_ sg13g2_buf_1
X_18899_ _11719_ _11641_ VPWR VGND _11720_ sg13g2_xnor2_1
X_18900_ _11637_ _11641_ _11656_ _11653_ VPWR VGND 
+ _11721_
+ sg13g2_a22oi_1
X_18901_ \atbs_core_0.dac_control_1.dac_counter_value[1]\ VPWR VGND _11722_ sg13g2_buf_1
X_18902_ _11722_ _11629_ _11440_ VPWR VGND _11723_ sg13g2_and3_1
X_18903_ _11631_ _11633_ _11723_ VPWR VGND _11724_ sg13g2_o21ai_1
X_18904_ _11722_ _11630_ _11385_ VPWR VGND _11725_ sg13g2_nor3_1
X_18905_ _11631_ _11633_ _11725_ VPWR VGND _11726_ sg13g2_o21ai_1
X_18906_ _08065_ _08267_ _08270_ _08044_ _11369_ VPWR 
+ VGND
+ _11727_ sg13g2_a221oi_1
X_18907_ _11724_ _11726_ _11727_ VPWR VGND _11728_ sg13g2_mux2_1
X_18908_ _11728_ VPWR VGND _11729_ sg13g2_buf_1
X_18909_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ VPWR VGND _11730_ sg13g2_buf_1
X_18910_ _11730_ _11661_ VPWR VGND _11731_ sg13g2_xnor2_1
X_18911_ _11642_ _11720_ _11721_ _11729_ _11731_ VPWR 
+ VGND
+ _11732_ sg13g2_a221oi_1
X_18912_ _11732_ VPWR VGND _11733_ sg13g2_buf_2
X_18913_ \atbs_core_0.dac_control_1.dac_counter_value[4]\ VPWR VGND _11734_ sg13g2_buf_1
X_18914_ _11734_ VPWR VGND _11735_ sg13g2_inv_1
X_18915_ _11673_ _11677_ VPWR VGND _11736_ sg13g2_nand2_1
X_18916_ _11735_ _11736_ VPWR VGND _11737_ sg13g2_nor2_1
X_18917_ _11718_ _11733_ _11737_ VPWR VGND _11738_ sg13g2_o21ai_1
X_18918_ _11738_ VPWR VGND _11739_ sg13g2_buf_1
X_18919_ _11673_ _11677_ VPWR VGND _11740_ sg13g2_and2_1
X_18920_ _11734_ _11740_ VPWR VGND _11741_ sg13g2_nor2_1
X_18921_ _11735_ _11662_ _11661_ VPWR VGND _11742_ sg13g2_nand3_1
X_18922_ _00098_ _11742_ _11740_ VPWR VGND _11743_ sg13g2_a21oi_1
X_18923_ _11733_ _11741_ _11669_ _11666_ _11743_ VPWR 
+ VGND
+ _11744_ sg13g2_a221oi_1
X_18924_ _11683_ _11685_ VPWR VGND _11745_ sg13g2_nor2_1
X_18925_ _11666_ _11669_ VPWR VGND _11746_ sg13g2_or2_1
X_18926_ _11745_ _11746_ VPWR VGND _11747_ sg13g2_nand2b_1
X_18927_ _11739_ _11744_ _11747_ VPWR VGND _11748_ sg13g2_a21oi_2
X_18928_ _11683_ _11685_ VPWR VGND _11749_ sg13g2_nand2_1
X_18929_ _11749_ VPWR VGND _11750_ sg13g2_inv_1
X_18930_ \atbs_core_0.dac_control_1.dac_counter_value[7]\ VPWR VGND _11751_ sg13g2_buf_1
X_18931_ _00099_ VPWR VGND _11752_ sg13g2_inv_1
X_18932_ _07936_ _11649_ _07843_ VPWR VGND _11753_ sg13g2_a21oi_1
X_18933_ _11751_ _11752_ _11753_ VPWR VGND _11754_ sg13g2_nand3_1
X_18934_ _11748_ _11750_ _11754_ VPWR VGND _11755_ sg13g2_or3_1
X_18935_ _11751_ _00099_ _11652_ VPWR VGND _11756_ sg13g2_nor3_1
X_18936_ _11748_ _11750_ _11756_ VPWR VGND _11757_ sg13g2_o21ai_1
X_18937_ _11707_ _07843_ VPWR VGND _11758_ sg13g2_nand2_1
X_18938_ _11755_ _11757_ _11758_ VPWR VGND _11759_ sg13g2_nand3_1
X_18939_ _11759_ VPWR VGND _11760_ sg13g2_buf_2
X_18940_ _11635_ _11715_ _11760_ VPWR VGND _11761_ sg13g2_a21oi_1
X_18941_ _11755_ _11757_ _11715_ VPWR VGND _11762_ sg13g2_nand3_1
X_18942_ _11762_ VPWR VGND _11763_ sg13g2_buf_2
X_18943_ _11763_ _11630_ _11647_ VPWR VGND _11764_ sg13g2_nand3b_1
X_18944_ _11630_ _11761_ _11764_ VPWR VGND _00566_ sg13g2_o21ai_1
X_18945_ _11722_ _11648_ VPWR VGND _11765_ sg13g2_xor2_1
X_18946_ _00097_ _11692_ VPWR VGND _11766_ sg13g2_xnor2_1
X_18947_ _11765_ _11766_ _11652_ VPWR VGND _11767_ sg13g2_mux2_1
X_18948_ _11689_ _11767_ VPWR VGND _11768_ sg13g2_xnor2_1
X_18949_ _11722_ _11760_ VPWR VGND _11769_ sg13g2_nand2_1
X_18950_ _11763_ _11768_ _11769_ VPWR VGND _00567_ sg13g2_o21ai_1
X_18951_ _11753_ VPWR VGND _11770_ sg13g2_buf_1
X_18952_ _00097_ _11689_ _11729_ VPWR VGND _11771_ sg13g2_o21ai_1
X_18953_ _11719_ _11771_ VPWR VGND _11772_ sg13g2_xor2_1
X_18954_ _11689_ _11692_ VPWR VGND _11773_ sg13g2_nand2_1
X_18955_ _11636_ _11694_ _11773_ VPWR VGND _11774_ sg13g2_nand3_1
X_18956_ _11694_ _11773_ _11636_ VPWR VGND _11775_ sg13g2_a21o_1
X_18957_ _11774_ _11775_ _11770_ VPWR VGND _11776_ sg13g2_a21oi_1
X_18958_ _11770_ _11772_ _11776_ VPWR VGND _11777_ sg13g2_a21oi_1
X_18959_ _11644_ _11777_ VPWR VGND _11778_ sg13g2_xnor2_1
X_18960_ _11719_ _11760_ VPWR VGND _11779_ sg13g2_nand2_1
X_18961_ _11763_ _11778_ _11779_ VPWR VGND _00568_ sg13g2_o21ai_1
X_18962_ _11642_ _11720_ _11721_ _11729_ VPWR VGND 
+ _11780_
+ sg13g2_a22oi_1
X_18963_ _11730_ _11780_ VPWR VGND _11781_ sg13g2_xnor2_1
X_18964_ _11662_ _11696_ VPWR VGND _11782_ sg13g2_xnor2_1
X_18965_ _11770_ _11782_ VPWR VGND _11783_ sg13g2_nor2_1
X_18966_ _11770_ _11781_ _11783_ VPWR VGND _11784_ sg13g2_a21oi_1
X_18967_ _11661_ _11784_ VPWR VGND _11785_ sg13g2_xnor2_1
X_18968_ _11730_ _11760_ VPWR VGND _11786_ sg13g2_nand2_1
X_18969_ _11763_ _11785_ _11786_ VPWR VGND _00569_ sg13g2_o21ai_1
X_18970_ _11718_ _11733_ VPWR VGND _11787_ sg13g2_nor2_1
X_18971_ _11735_ _11787_ VPWR VGND _11788_ sg13g2_xnor2_1
X_18972_ _11637_ _11644_ _11662_ VPWR VGND _11789_ sg13g2_o21ai_1
X_18973_ _11636_ _11641_ _11661_ VPWR VGND _11790_ sg13g2_a21o_1
X_18974_ _11694_ _11695_ _11789_ _11790_ VPWR VGND 
+ _11791_
+ sg13g2_a22oi_1
X_18975_ _11791_ _11663_ VPWR VGND _11792_ sg13g2_nand2b_1
X_18976_ _11678_ _11792_ VPWR VGND _11793_ sg13g2_xnor2_1
X_18977_ _11770_ _11793_ VPWR VGND _11794_ sg13g2_nor2_1
X_18978_ _11770_ _11788_ _11794_ VPWR VGND _11795_ sg13g2_a21oi_1
X_18979_ _11736_ _11795_ VPWR VGND _11796_ sg13g2_xnor2_1
X_18980_ _11734_ _11760_ VPWR VGND _11797_ sg13g2_nand2_1
X_18981_ _11763_ _11796_ _11797_ VPWR VGND _00570_ sg13g2_o21ai_1
X_18982_ _11770_ _11739_ VPWR VGND _11798_ sg13g2_nand2_1
X_18983_ _11678_ _11792_ _11652_ VPWR VGND _11799_ sg13g2_o21ai_1
X_18984_ _11678_ _11652_ VPWR VGND _11800_ sg13g2_nor2_1
X_18985_ _11718_ _11733_ _11735_ VPWR VGND _11801_ sg13g2_o21ai_1
X_18986_ _00098_ _11753_ VPWR VGND _11802_ sg13g2_nor2_1
X_18987_ _11800_ _11801_ _11802_ _11792_ VPWR VGND 
+ _11803_
+ sg13g2_a22oi_1
X_18988_ _11798_ _11799_ _11803_ _11736_ VPWR VGND 
+ _11804_
+ sg13g2_a22oi_1
X_18989_ _11669_ _11804_ VPWR VGND _11805_ sg13g2_xor2_1
X_18990_ _11715_ _11805_ _11760_ VPWR VGND _11806_ sg13g2_a21o_1
X_18991_ _11666_ _11763_ _11805_ VPWR VGND _11807_ sg13g2_nor3_1
X_18992_ _11666_ _11806_ _11807_ VPWR VGND _00571_ sg13g2_a21o_1
X_18993_ _11698_ _11710_ VPWR VGND _11808_ sg13g2_nand2_1
X_18994_ _00036_ _11652_ VPWR VGND _11809_ sg13g2_nand2b_1
X_18995_ _11770_ _11746_ VPWR VGND _11810_ sg13g2_nand2_1
X_18996_ _11739_ _11744_ _11810_ VPWR VGND _11811_ sg13g2_a21o_1
X_18997_ _11808_ _11809_ _11811_ VPWR VGND _11812_ sg13g2_o21ai_1
X_18998_ _11770_ _11703_ _11705_ VPWR VGND _11813_ sg13g2_nor3_1
X_18999_ _11683_ _11685_ _11701_ VPWR VGND _11814_ sg13g2_nand3b_1
X_19000_ _11683_ _11700_ VPWR VGND _11815_ sg13g2_nand2_1
X_19001_ _11698_ _11813_ _11814_ _11815_ VPWR VGND 
+ _11816_
+ sg13g2_a22oi_1
X_19002_ _11745_ _11812_ _11816_ _11811_ VPWR VGND 
+ _11817_
+ sg13g2_a22oi_1
X_19003_ _11707_ \atbs_core_0.dac_control_1.dac_init_value[6]\ VPWR VGND _11818_ sg13g2_nor2_1
X_19004_ _11707_ _11817_ _11818_ VPWR VGND _11819_ sg13g2_a21o_1
X_19005_ _11707_ _11685_ _11812_ VPWR VGND _11820_ sg13g2_and3_1
X_19006_ _11760_ _11820_ _11683_ VPWR VGND _11821_ sg13g2_o21ai_1
X_19007_ _11760_ _11819_ _11821_ VPWR VGND _00572_ sg13g2_o21ai_1
X_19008_ _11748_ _11749_ VPWR VGND _11822_ sg13g2_nand2b_1
X_19009_ _11751_ _11752_ _11652_ VPWR VGND _11823_ sg13g2_nor3_1
X_19010_ _11700_ _11808_ VPWR VGND _11824_ sg13g2_nand2_1
X_19011_ _11700_ _11808_ _11683_ VPWR VGND _11825_ sg13g2_o21ai_1
X_19012_ _11824_ _11825_ _11809_ VPWR VGND _11826_ sg13g2_a21oi_1
X_19013_ _11822_ _11823_ _11826_ VPWR VGND _11827_ sg13g2_a21oi_1
X_19014_ _11752_ _11707_ _11770_ VPWR VGND _11828_ sg13g2_o21ai_1
X_19015_ _11822_ _11828_ _11758_ VPWR VGND _11829_ sg13g2_o21ai_1
X_19016_ _11751_ _11829_ VPWR VGND _11830_ sg13g2_nand2_1
X_19017_ _11708_ _11827_ _11830_ VPWR VGND _00573_ sg13g2_o21ai_1
X_19018_ \atbs_core_0.dac_control_1.n2091_q[1]\ \atbs_core_0.dac_control_1.n2091_q[0]\ VPWR VGND _11831_ sg13g2_nand2_1
X_19019_ _00059_ _11831_ VPWR VGND _11832_ sg13g2_or2_1
X_19020_ _11707_ VPWR VGND _11833_ sg13g2_inv_1
X_19021_ \atbs_core_0.dac_control_1.n1981_o\ _11833_ _07843_ VPWR VGND _11834_ sg13g2_a21oi_1
X_19022_ \atbs_core_0.dac_control_1.dac_change_in_progress\ _11832_ _11834_ VPWR VGND _00574_ sg13g2_a21o_1
X_19023_ dac_lower_o[0] VPWR VGND _11835_ sg13g2_inv_1
X_19024_ _07843_ _11736_ _11669_ _11685_ VPWR VGND 
+ _11836_
+ sg13g2_nor4_1
X_19025_ _11717_ _11836_ VPWR VGND _11837_ sg13g2_and2_1
X_19026_ _11837_ VPWR VGND _11838_ sg13g2_buf_1
X_19027_ _11635_ _11641_ _11656_ VPWR VGND _11839_ sg13g2_nor3_1
X_19028_ _11835_ _07843_ _11838_ _11839_ VPWR VGND 
+ _00575_
+ sg13g2_a22oi_1
X_19029_ dac_lower_o[1] VPWR VGND _11840_ sg13g2_inv_1
X_19030_ _11635_ _11689_ VPWR VGND _11841_ sg13g2_xnor2_1
X_19031_ _11641_ _11841_ VPWR VGND _11842_ sg13g2_nor2_1
X_19032_ _11840_ _07843_ _11838_ _11842_ VPWR VGND 
+ _00576_
+ sg13g2_a22oi_1
X_19033_ dac_lower_o[2] VPWR VGND _11843_ sg13g2_inv_1
X_19034_ _11635_ _11641_ _11689_ VPWR VGND _11844_ sg13g2_nand3_1
X_19035_ _11641_ _11841_ _11844_ VPWR VGND _11845_ sg13g2_o21ai_1
X_19036_ _11843_ _07843_ _11838_ _11845_ VPWR VGND 
+ _00577_
+ sg13g2_a22oi_1
X_19037_ dac_lower_o[3] VPWR VGND _11846_ sg13g2_inv_1
X_19038_ _11661_ _11845_ VPWR VGND _11847_ sg13g2_nor2_1
X_19039_ _11641_ _11656_ VPWR VGND _11848_ sg13g2_nor2_1
X_19040_ _11635_ _11848_ _11717_ VPWR VGND _11849_ sg13g2_a21oi_1
X_19041_ _11847_ _11849_ VPWR VGND _11850_ sg13g2_nor2_1
X_19042_ _11846_ _07843_ _11836_ _11850_ VPWR VGND 
+ _00578_
+ sg13g2_a22oi_1
X_19043_ \atbs_core_0.debouncer_0.n1511_q[1]\ VPWR VGND _11851_ sg13g2_buf_1
X_19044_ \atbs_core_0.debouncer_0.n1511_q[0]\ VPWR VGND _11852_ sg13g2_buf_1
X_19045_ \atbs_core_0.debouncer_0.counter_value[10]\ VPWR VGND _11853_ sg13g2_inv_1
X_19046_ \atbs_core_0.debouncer_0.counter_value[3]\ VPWR VGND _11854_ sg13g2_inv_1
X_19047_ \atbs_core_0.debouncer_0.counter_value[0]\ VPWR VGND _11855_ sg13g2_buf_1
X_19048_ \atbs_core_0.debouncer_0.counter_value[1]\ _11855_ \atbs_core_0.debouncer_0.counter_value[2]\ VPWR VGND _11856_ sg13g2_nand3_1
X_19049_ _11854_ _11856_ VPWR VGND _11857_ sg13g2_nor2_1
X_19050_ \atbs_core_0.debouncer_0.counter_value[5]\ \atbs_core_0.debouncer_0.counter_value[4]\ _11857_ VPWR VGND _11858_ sg13g2_and3_1
X_19051_ _11858_ VPWR VGND _11859_ sg13g2_buf_1
X_19052_ \atbs_core_0.debouncer_0.counter_value[7]\ \atbs_core_0.debouncer_0.counter_value[6]\ _11859_ VPWR VGND _11860_ sg13g2_and3_1
X_19053_ _11860_ VPWR VGND _11861_ sg13g2_buf_1
X_19054_ \atbs_core_0.debouncer_0.counter_value[9]\ \atbs_core_0.debouncer_0.counter_value[8]\ _11861_ VPWR VGND _11862_ sg13g2_nand3_1
X_19055_ _11853_ _11862_ VPWR VGND _11863_ sg13g2_nor2_1
X_19056_ \atbs_core_0.debouncer_0.counter_value[11]\ _11863_ VPWR VGND _11864_ sg13g2_and2_1
X_19057_ _11864_ VPWR VGND _11865_ sg13g2_buf_1
X_19058_ \atbs_core_0.debouncer_0.counter_value[13]\ \atbs_core_0.debouncer_0.counter_value[12]\ _11865_ VPWR VGND _11866_ sg13g2_and3_1
X_19059_ _11866_ VPWR VGND _11867_ sg13g2_buf_1
X_19060_ \atbs_core_0.debouncer_0.counter_value[14]\ \atbs_core_0.debouncer_0.counter_value[15]\ _11867_ VPWR VGND _11868_ sg13g2_nand3_1
X_19061_ _11868_ VPWR VGND _11869_ sg13g2_buf_1
X_19062_ \atbs_core_0.debouncer_0.bouncing_sync_d\ VPWR VGND _11870_ sg13g2_buf_1
X_19063_ _11870_ VPWR VGND _11871_ sg13g2_inv_1
X_19064_ _11852_ \atbs_core_0.debouncer_0.bouncing_sync\ _11871_ VPWR VGND _11872_ sg13g2_nor3_1
X_19065_ _11852_ _11869_ _11872_ VPWR VGND _11873_ sg13g2_a21oi_1
X_19066_ _11851_ _11873_ VPWR VGND _00579_ sg13g2_nor2_1
X_19067_ \atbs_core_0.debouncer_0.bouncing_sync\ VPWR VGND _11874_ sg13g2_inv_1
X_19068_ _11851_ _11874_ _11870_ VPWR VGND _11875_ sg13g2_nor3_1
X_19069_ _11851_ _11869_ _11875_ VPWR VGND _11876_ sg13g2_a21oi_1
X_19070_ _11852_ _11876_ VPWR VGND _00580_ sg13g2_nor2_1
X_19071_ _11852_ _11851_ VPWR VGND _11877_ sg13g2_xnor2_1
X_19072_ _11869_ _11877_ VPWR VGND _11878_ sg13g2_nor2_1
X_19073_ \atbs_core_0.debouncer_0.debounced\ _11870_ _11878_ VPWR VGND _00581_ sg13g2_mux2_1
X_19074_ \atbs_core_0.debouncer_1.n1511_q[1]\ VPWR VGND _11879_ sg13g2_buf_1
X_19075_ \atbs_core_0.debouncer_1.n1511_q[0]\ VPWR VGND _11880_ sg13g2_buf_1
X_19076_ \atbs_core_0.debouncer_1.counter_value[10]\ VPWR VGND _11881_ sg13g2_inv_1
X_19077_ \atbs_core_0.debouncer_1.counter_value[3]\ VPWR VGND _11882_ sg13g2_inv_1
X_19078_ \atbs_core_0.debouncer_1.counter_value[0]\ VPWR VGND _11883_ sg13g2_buf_1
X_19079_ \atbs_core_0.debouncer_1.counter_value[1]\ _11883_ \atbs_core_0.debouncer_1.counter_value[2]\ VPWR VGND _11884_ sg13g2_nand3_1
X_19080_ _11882_ _11884_ VPWR VGND _11885_ sg13g2_nor2_1
X_19081_ \atbs_core_0.debouncer_1.counter_value[5]\ \atbs_core_0.debouncer_1.counter_value[4]\ _11885_ VPWR VGND _11886_ sg13g2_and3_1
X_19082_ _11886_ VPWR VGND _11887_ sg13g2_buf_1
X_19083_ \atbs_core_0.debouncer_1.counter_value[7]\ \atbs_core_0.debouncer_1.counter_value[6]\ _11887_ VPWR VGND _11888_ sg13g2_and3_1
X_19084_ _11888_ VPWR VGND _11889_ sg13g2_buf_1
X_19085_ \atbs_core_0.debouncer_1.counter_value[9]\ \atbs_core_0.debouncer_1.counter_value[8]\ _11889_ VPWR VGND _11890_ sg13g2_nand3_1
X_19086_ _11881_ _11890_ VPWR VGND _11891_ sg13g2_nor2_1
X_19087_ \atbs_core_0.debouncer_1.counter_value[11]\ _11891_ VPWR VGND _11892_ sg13g2_and2_1
X_19088_ _11892_ VPWR VGND _11893_ sg13g2_buf_1
X_19089_ \atbs_core_0.debouncer_1.counter_value[13]\ \atbs_core_0.debouncer_1.counter_value[12]\ _11893_ VPWR VGND _11894_ sg13g2_and3_1
X_19090_ _11894_ VPWR VGND _11895_ sg13g2_buf_1
X_19091_ \atbs_core_0.debouncer_1.counter_value[14]\ \atbs_core_0.debouncer_1.counter_value[15]\ _11895_ VPWR VGND _11896_ sg13g2_nand3_1
X_19092_ _11896_ VPWR VGND _11897_ sg13g2_buf_1
X_19093_ \atbs_core_0.debouncer_1.bouncing_sync_d\ VPWR VGND _11898_ sg13g2_buf_1
X_19094_ _11898_ VPWR VGND _11899_ sg13g2_inv_1
X_19095_ _11880_ \atbs_core_0.debouncer_1.bouncing_sync\ _11899_ VPWR VGND _11900_ sg13g2_nor3_1
X_19096_ _11880_ _11897_ _11900_ VPWR VGND _11901_ sg13g2_a21oi_1
X_19097_ _11879_ _11901_ VPWR VGND _00582_ sg13g2_nor2_1
X_19098_ \atbs_core_0.debouncer_1.bouncing_sync\ VPWR VGND _11902_ sg13g2_inv_1
X_19099_ _11879_ _11902_ _11898_ VPWR VGND _11903_ sg13g2_nor3_1
X_19100_ _11879_ _11897_ _11903_ VPWR VGND _11904_ sg13g2_a21oi_1
X_19101_ _11880_ _11904_ VPWR VGND _00583_ sg13g2_nor2_1
X_19102_ _11880_ _11879_ VPWR VGND _11905_ sg13g2_xnor2_1
X_19103_ _11897_ _11905_ VPWR VGND _11906_ sg13g2_nor2_1
X_19104_ _07710_ _11898_ _11906_ VPWR VGND _00584_ sg13g2_mux2_1
X_19105_ \atbs_core_0.debouncer_2.n1511_q[1]\ VPWR VGND _11907_ sg13g2_buf_1
X_19106_ \atbs_core_0.debouncer_2.n1511_q[0]\ VPWR VGND _11908_ sg13g2_buf_1
X_19107_ \atbs_core_0.debouncer_2.counter_value[10]\ VPWR VGND _11909_ sg13g2_inv_1
X_19108_ \atbs_core_0.debouncer_2.counter_value[3]\ VPWR VGND _11910_ sg13g2_inv_1
X_19109_ \atbs_core_0.debouncer_2.counter_value[0]\ VPWR VGND _11911_ sg13g2_buf_1
X_19110_ \atbs_core_0.debouncer_2.counter_value[1]\ _11911_ \atbs_core_0.debouncer_2.counter_value[2]\ VPWR VGND _11912_ sg13g2_nand3_1
X_19111_ _11910_ _11912_ VPWR VGND _11913_ sg13g2_nor2_1
X_19112_ \atbs_core_0.debouncer_2.counter_value[5]\ \atbs_core_0.debouncer_2.counter_value[4]\ _11913_ VPWR VGND _11914_ sg13g2_and3_1
X_19113_ _11914_ VPWR VGND _11915_ sg13g2_buf_1
X_19114_ \atbs_core_0.debouncer_2.counter_value[7]\ \atbs_core_0.debouncer_2.counter_value[6]\ _11915_ VPWR VGND _11916_ sg13g2_and3_1
X_19115_ _11916_ VPWR VGND _11917_ sg13g2_buf_1
X_19116_ \atbs_core_0.debouncer_2.counter_value[9]\ \atbs_core_0.debouncer_2.counter_value[8]\ _11917_ VPWR VGND _11918_ sg13g2_nand3_1
X_19117_ _11909_ _11918_ VPWR VGND _11919_ sg13g2_nor2_1
X_19118_ \atbs_core_0.debouncer_2.counter_value[11]\ _11919_ VPWR VGND _11920_ sg13g2_and2_1
X_19119_ _11920_ VPWR VGND _11921_ sg13g2_buf_1
X_19120_ \atbs_core_0.debouncer_2.counter_value[13]\ \atbs_core_0.debouncer_2.counter_value[12]\ _11921_ VPWR VGND _11922_ sg13g2_and3_1
X_19121_ _11922_ VPWR VGND _11923_ sg13g2_buf_1
X_19122_ \atbs_core_0.debouncer_2.counter_value[14]\ \atbs_core_0.debouncer_2.counter_value[15]\ _11923_ VPWR VGND _11924_ sg13g2_nand3_1
X_19123_ _11924_ VPWR VGND _11925_ sg13g2_buf_1
X_19124_ \atbs_core_0.debouncer_2.bouncing_sync_d\ VPWR VGND _11926_ sg13g2_buf_1
X_19125_ _11926_ VPWR VGND _11927_ sg13g2_inv_1
X_19126_ _11908_ \atbs_core_0.debouncer_2.bouncing_sync\ _11927_ VPWR VGND _11928_ sg13g2_nor3_1
X_19127_ _11908_ _11925_ _11928_ VPWR VGND _11929_ sg13g2_a21oi_1
X_19128_ _11907_ _11929_ VPWR VGND _00585_ sg13g2_nor2_1
X_19129_ \atbs_core_0.debouncer_2.bouncing_sync\ VPWR VGND _11930_ sg13g2_inv_1
X_19130_ _11907_ _11930_ _11926_ VPWR VGND _11931_ sg13g2_nor3_1
X_19131_ _11907_ _11925_ _11931_ VPWR VGND _11932_ sg13g2_a21oi_1
X_19132_ _11908_ _11932_ VPWR VGND _00586_ sg13g2_nor2_1
X_19133_ _11908_ _11907_ VPWR VGND _11933_ sg13g2_xnor2_1
X_19134_ _11925_ _11933_ VPWR VGND _11934_ sg13g2_nor2_1
X_19135_ _07653_ _11926_ _11934_ VPWR VGND _00587_ sg13g2_mux2_1
X_19136_ \atbs_core_0.debouncer_3.n1511_q[1]\ VPWR VGND _11935_ sg13g2_buf_1
X_19137_ \atbs_core_0.debouncer_3.n1511_q[0]\ VPWR VGND _11936_ sg13g2_buf_1
X_19138_ \atbs_core_0.debouncer_3.counter_value[14]\ VPWR VGND _11937_ sg13g2_inv_1
X_19139_ \atbs_core_0.debouncer_3.counter_value[11]\ VPWR VGND _11938_ sg13g2_inv_1
X_19140_ \atbs_core_0.debouncer_3.counter_value[8]\ VPWR VGND _11939_ sg13g2_inv_1
X_19141_ \atbs_core_0.debouncer_3.counter_value[3]\ VPWR VGND _11940_ sg13g2_inv_1
X_19142_ \atbs_core_0.debouncer_3.counter_value[0]\ VPWR VGND _11941_ sg13g2_buf_1
X_19143_ \atbs_core_0.debouncer_3.counter_value[1]\ _11941_ \atbs_core_0.debouncer_3.counter_value[2]\ VPWR VGND _11942_ sg13g2_nand3_1
X_19144_ _11940_ _11942_ VPWR VGND _11943_ sg13g2_nor2_1
X_19145_ \atbs_core_0.debouncer_3.counter_value[5]\ \atbs_core_0.debouncer_3.counter_value[4]\ _11943_ VPWR VGND _11944_ sg13g2_and3_1
X_19146_ _11944_ VPWR VGND _11945_ sg13g2_buf_1
X_19147_ \atbs_core_0.debouncer_3.counter_value[7]\ \atbs_core_0.debouncer_3.counter_value[6]\ _11945_ VPWR VGND _11946_ sg13g2_nand3_1
X_19148_ _11939_ _11946_ VPWR VGND _11947_ sg13g2_nor2_1
X_19149_ \atbs_core_0.debouncer_3.counter_value[9]\ \atbs_core_0.debouncer_3.counter_value[10]\ _11947_ VPWR VGND _11948_ sg13g2_nand3_1
X_19150_ _11938_ _11948_ VPWR VGND _11949_ sg13g2_nor2_1
X_19151_ \atbs_core_0.debouncer_3.counter_value[13]\ \atbs_core_0.debouncer_3.counter_value[12]\ _11949_ VPWR VGND _11950_ sg13g2_nand3_1
X_19152_ _11937_ _11950_ VPWR VGND _11951_ sg13g2_nor2_1
X_19153_ \atbs_core_0.debouncer_3.counter_value[15]\ _11951_ VPWR VGND _11952_ sg13g2_nand2_1
X_19154_ \atbs_core_0.debouncer_3.bouncing_sync_d\ VPWR VGND _11953_ sg13g2_buf_1
X_19155_ _11953_ VPWR VGND _11954_ sg13g2_inv_1
X_19156_ _11936_ \atbs_core_0.debouncer_3.bouncing_sync\ _11954_ VPWR VGND _11955_ sg13g2_nor3_1
X_19157_ _11936_ _11952_ _11955_ VPWR VGND _11956_ sg13g2_a21oi_1
X_19158_ _11935_ _11956_ VPWR VGND _00588_ sg13g2_nor2_1
X_19159_ \atbs_core_0.debouncer_3.bouncing_sync\ VPWR VGND _11957_ sg13g2_inv_1
X_19160_ _11935_ _11957_ _11953_ VPWR VGND _11958_ sg13g2_nor3_1
X_19161_ _11935_ _11952_ _11958_ VPWR VGND _11959_ sg13g2_a21oi_1
X_19162_ _11936_ _11959_ VPWR VGND _00589_ sg13g2_nor2_1
X_19163_ _11936_ _11935_ VPWR VGND _11960_ sg13g2_xnor2_1
X_19164_ _11952_ _11960_ VPWR VGND _11961_ sg13g2_nor2_1
X_19165_ \atbs_core_0.debouncer_3.debounced\ _11953_ _11961_ VPWR VGND _00590_ sg13g2_mux2_1
X_19166_ \atbs_core_0.debouncer_4.n1511_q[1]\ VPWR VGND _11962_ sg13g2_buf_1
X_19167_ \atbs_core_0.debouncer_4.n1511_q[0]\ VPWR VGND _11963_ sg13g2_buf_1
X_19168_ \atbs_core_0.debouncer_4.counter_value[14]\ VPWR VGND _11964_ sg13g2_inv_1
X_19169_ \atbs_core_0.debouncer_4.counter_value[11]\ VPWR VGND _11965_ sg13g2_inv_1
X_19170_ \atbs_core_0.debouncer_4.counter_value[8]\ VPWR VGND _11966_ sg13g2_inv_1
X_19171_ \atbs_core_0.debouncer_4.counter_value[3]\ VPWR VGND _11967_ sg13g2_inv_1
X_19172_ \atbs_core_0.debouncer_4.counter_value[0]\ VPWR VGND _11968_ sg13g2_buf_1
X_19173_ \atbs_core_0.debouncer_4.counter_value[1]\ _11968_ \atbs_core_0.debouncer_4.counter_value[2]\ VPWR VGND _11969_ sg13g2_nand3_1
X_19174_ _11967_ _11969_ VPWR VGND _11970_ sg13g2_nor2_1
X_19175_ \atbs_core_0.debouncer_4.counter_value[5]\ \atbs_core_0.debouncer_4.counter_value[4]\ _11970_ VPWR VGND _11971_ sg13g2_and3_1
X_19176_ _11971_ VPWR VGND _11972_ sg13g2_buf_1
X_19177_ \atbs_core_0.debouncer_4.counter_value[7]\ \atbs_core_0.debouncer_4.counter_value[6]\ _11972_ VPWR VGND _11973_ sg13g2_nand3_1
X_19178_ _11966_ _11973_ VPWR VGND _11974_ sg13g2_nor2_1
X_19179_ \atbs_core_0.debouncer_4.counter_value[9]\ \atbs_core_0.debouncer_4.counter_value[10]\ _11974_ VPWR VGND _11975_ sg13g2_nand3_1
X_19180_ _11965_ _11975_ VPWR VGND _11976_ sg13g2_nor2_1
X_19181_ \atbs_core_0.debouncer_4.counter_value[13]\ \atbs_core_0.debouncer_4.counter_value[12]\ _11976_ VPWR VGND _11977_ sg13g2_nand3_1
X_19182_ _11964_ _11977_ VPWR VGND _11978_ sg13g2_nor2_1
X_19183_ \atbs_core_0.debouncer_4.counter_value[15]\ _11978_ VPWR VGND _11979_ sg13g2_nand2_1
X_19184_ \atbs_core_0.debouncer_4.bouncing_sync_d\ VPWR VGND _11980_ sg13g2_buf_1
X_19185_ _11980_ VPWR VGND _11981_ sg13g2_inv_1
X_19186_ \atbs_core_0.debouncer_4.bouncing_sync\ _11981_ _11963_ VPWR VGND _11982_ sg13g2_nor3_1
X_19187_ _11963_ _11979_ _11982_ VPWR VGND _11983_ sg13g2_a21oi_1
X_19188_ _11962_ _11983_ VPWR VGND _00591_ sg13g2_nor2_1
X_19189_ \atbs_core_0.debouncer_4.bouncing_sync\ VPWR VGND _11984_ sg13g2_inv_1
X_19190_ _11984_ _11980_ _11962_ VPWR VGND _11985_ sg13g2_nor3_1
X_19191_ _11962_ _11979_ _11985_ VPWR VGND _11986_ sg13g2_a21oi_1
X_19192_ _11963_ _11986_ VPWR VGND _00592_ sg13g2_nor2_1
X_19193_ _11963_ _11962_ VPWR VGND _11987_ sg13g2_xnor2_1
X_19194_ _11979_ _11987_ VPWR VGND _11988_ sg13g2_nor2_1
X_19195_ \atbs_core_0.debouncer_4.debounced\ _11980_ _11988_ VPWR VGND _00593_ sg13g2_mux2_1
X_19196_ \atbs_core_0.debouncer_5.n1511_q[1]\ VPWR VGND _11989_ sg13g2_buf_1
X_19197_ \atbs_core_0.debouncer_5.n1511_q[0]\ VPWR VGND _11990_ sg13g2_buf_1
X_19198_ \atbs_core_0.debouncer_5.counter_value[10]\ VPWR VGND _11991_ sg13g2_inv_1
X_19199_ \atbs_core_0.debouncer_5.counter_value[3]\ VPWR VGND _11992_ sg13g2_inv_1
X_19200_ \atbs_core_0.debouncer_5.counter_value[0]\ VPWR VGND _11993_ sg13g2_buf_1
X_19201_ \atbs_core_0.debouncer_5.counter_value[1]\ _11993_ \atbs_core_0.debouncer_5.counter_value[2]\ VPWR VGND _11994_ sg13g2_nand3_1
X_19202_ _11992_ _11994_ VPWR VGND _11995_ sg13g2_nor2_1
X_19203_ \atbs_core_0.debouncer_5.counter_value[5]\ \atbs_core_0.debouncer_5.counter_value[4]\ _11995_ VPWR VGND _11996_ sg13g2_and3_1
X_19204_ _11996_ VPWR VGND _11997_ sg13g2_buf_1
X_19205_ \atbs_core_0.debouncer_5.counter_value[7]\ \atbs_core_0.debouncer_5.counter_value[6]\ _11997_ VPWR VGND _11998_ sg13g2_and3_1
X_19206_ _11998_ VPWR VGND _11999_ sg13g2_buf_1
X_19207_ \atbs_core_0.debouncer_5.counter_value[9]\ \atbs_core_0.debouncer_5.counter_value[8]\ _11999_ VPWR VGND _12000_ sg13g2_nand3_1
X_19208_ _11991_ _12000_ VPWR VGND _12001_ sg13g2_nor2_1
X_19209_ \atbs_core_0.debouncer_5.counter_value[11]\ _12001_ VPWR VGND _12002_ sg13g2_and2_1
X_19210_ _12002_ VPWR VGND _12003_ sg13g2_buf_1
X_19211_ \atbs_core_0.debouncer_5.counter_value[13]\ \atbs_core_0.debouncer_5.counter_value[12]\ _12003_ VPWR VGND _12004_ sg13g2_and3_1
X_19212_ _12004_ VPWR VGND _12005_ sg13g2_buf_1
X_19213_ \atbs_core_0.debouncer_5.counter_value[14]\ \atbs_core_0.debouncer_5.counter_value[15]\ _12005_ VPWR VGND _12006_ sg13g2_nand3_1
X_19214_ _12006_ VPWR VGND _12007_ sg13g2_buf_1
X_19215_ \atbs_core_0.debouncer_5.bouncing_sync_d\ VPWR VGND _12008_ sg13g2_buf_1
X_19216_ _12008_ VPWR VGND _12009_ sg13g2_inv_1
X_19217_ _11990_ \atbs_core_0.debouncer_5.bouncing_sync\ _12009_ VPWR VGND _12010_ sg13g2_nor3_1
X_19218_ _11990_ _12007_ _12010_ VPWR VGND _12011_ sg13g2_a21oi_1
X_19219_ _11989_ _12011_ VPWR VGND _00594_ sg13g2_nor2_1
X_19220_ \atbs_core_0.debouncer_5.bouncing_sync\ VPWR VGND _12012_ sg13g2_inv_1
X_19221_ _11989_ _12012_ _12008_ VPWR VGND _12013_ sg13g2_nor3_1
X_19222_ _11989_ _12007_ _12013_ VPWR VGND _12014_ sg13g2_a21oi_1
X_19223_ _11990_ _12014_ VPWR VGND _00595_ sg13g2_nor2_1
X_19224_ _11989_ _11990_ VPWR VGND _12015_ sg13g2_xnor2_1
X_19225_ _12007_ _12015_ VPWR VGND _12016_ sg13g2_nor2_1
X_19226_ \atbs_core_0.debouncer_5.debounced\ _12008_ _12016_ VPWR VGND _00596_ sg13g2_mux2_1
X_19227_ \atbs_core_0.memory2uart_0.tx_strb_i\ VPWR VGND _12017_ sg13g2_buf_1
X_19228_ _12017_ VPWR VGND _12018_ sg13g2_inv_1
X_19229_ \atbs_core_0.memory2uart_0.read_strb_i\ VPWR VGND _12019_ sg13g2_buf_1
X_19230_ _12019_ VPWR VGND _12020_ sg13g2_inv_1
X_19231_ _12018_ \atbs_core_0.memory2uart_0.counter[1]\ _12020_ VPWR VGND \atbs_core_0.memory2uart_0.n2588_o\ sg13g2_o21ai_1
X_19232_ _12019_ VPWR VGND _12021_ sg13g2_buf_1
X_19233_ _12021_ VPWR VGND _12022_ sg13g2_buf_1
X_19234_ _12018_ \atbs_core_0.memory2uart_0.counter[1]\ VPWR VGND _12023_ sg13g2_nor2_1
X_19235_ _12023_ VPWR VGND _12024_ sg13g2_buf_1
X_19236_ _12024_ VPWR VGND _12025_ sg13g2_buf_1
X_19237_ _12024_ VPWR VGND _12026_ sg13g2_buf_1
X_19238_ _12026_ \atbs_core_0.uart_0.uart_tx_0.n3348_o\ VPWR VGND _12027_ sg13g2_nor2b_1
X_19239_ \atbs_core_0.memory2uart_0.n2574_o[0]\ _12025_ _12027_ VPWR VGND _12028_ sg13g2_a21oi_1
X_19240_ _12021_ VPWR VGND _12029_ sg13g2_buf_1
X_19241_ _12029_ \atbs_core_0.b_data[16]\ VPWR VGND _12030_ sg13g2_nand2_1
X_19242_ _12022_ _12028_ _12030_ VPWR VGND _00597_ sg13g2_o21ai_1
X_19243_ _12026_ \atbs_core_0.memory2uart_0.n2574_o[2]\ VPWR VGND _12031_ sg13g2_nor2b_1
X_19244_ \atbs_core_0.memory2uart_0.n2574_o[10]\ _12025_ _12031_ VPWR VGND _12032_ sg13g2_a21oi_1
X_19245_ _12029_ \atbs_core_0.b_data[10]\ VPWR VGND _12033_ sg13g2_nand2_1
X_19246_ _12022_ _12032_ _12033_ VPWR VGND _00598_ sg13g2_o21ai_1
X_19247_ _12024_ VPWR VGND _12034_ sg13g2_buf_1
X_19248_ _12026_ \atbs_core_0.memory2uart_0.n2574_o[3]\ VPWR VGND _12035_ sg13g2_nor2b_1
X_19249_ \atbs_core_0.memory2uart_0.n2574_o[11]\ _12034_ _12035_ VPWR VGND _12036_ sg13g2_a21oi_1
X_19250_ _12021_ \atbs_core_0.b_data[11]\ VPWR VGND _12037_ sg13g2_nand2_1
X_19251_ _12022_ _12036_ _12037_ VPWR VGND _00599_ sg13g2_o21ai_1
X_19252_ _12026_ \atbs_core_0.memory2uart_0.n2574_o[4]\ VPWR VGND _12038_ sg13g2_nor2b_1
X_19253_ \atbs_core_0.memory2uart_0.n2574_o[12]\ _12034_ _12038_ VPWR VGND _12039_ sg13g2_a21oi_1
X_19254_ _12021_ \atbs_core_0.b_data[12]\ VPWR VGND _12040_ sg13g2_nand2_1
X_19255_ _12022_ _12039_ _12040_ VPWR VGND _00600_ sg13g2_o21ai_1
X_19256_ _12026_ \atbs_core_0.memory2uart_0.n2574_o[5]\ VPWR VGND _12041_ sg13g2_nor2b_1
X_19257_ \atbs_core_0.memory2uart_0.n2574_o[13]\ _12034_ _12041_ VPWR VGND _12042_ sg13g2_a21oi_1
X_19258_ _12021_ \atbs_core_0.b_data[13]\ VPWR VGND _12043_ sg13g2_nand2_1
X_19259_ _12022_ _12042_ _12043_ VPWR VGND _00601_ sg13g2_o21ai_1
X_19260_ _12026_ \atbs_core_0.memory2uart_0.n2574_o[6]\ VPWR VGND _12044_ sg13g2_nor2b_1
X_19261_ \atbs_core_0.memory2uart_0.n2574_o[14]\ _12034_ _12044_ VPWR VGND _12045_ sg13g2_a21oi_1
X_19262_ _12021_ \atbs_core_0.b_data[14]\ VPWR VGND _12046_ sg13g2_nand2_1
X_19263_ _12022_ _12045_ _12046_ VPWR VGND _00602_ sg13g2_o21ai_1
X_19264_ _12024_ \atbs_core_0.memory2uart_0.n2574_o[7]\ VPWR VGND _12047_ sg13g2_nor2b_1
X_19265_ \atbs_core_0.memory2uart_0.n2574_o[15]\ _12034_ _12047_ VPWR VGND _12048_ sg13g2_a21oi_1
X_19266_ _12021_ \atbs_core_0.b_data[15]\ VPWR VGND _12049_ sg13g2_nand2_1
X_19267_ _12022_ _12048_ _12049_ VPWR VGND _00603_ sg13g2_o21ai_1
X_19268_ \atbs_core_0.memory2uart_0.n2574_o[8]\ \atbs_core_0.b_data[0]\ _12029_ VPWR VGND _00604_ sg13g2_mux2_1
X_19269_ \atbs_core_0.memory2uart_0.n2574_o[9]\ \atbs_core_0.b_data[1]\ _12029_ VPWR VGND _00605_ sg13g2_mux2_1
X_19270_ \atbs_core_0.memory2uart_0.n2574_o[10]\ \atbs_core_0.b_data[2]\ _12029_ VPWR VGND _00606_ sg13g2_mux2_1
X_19271_ \atbs_core_0.memory2uart_0.n2574_o[11]\ \atbs_core_0.b_data[3]\ _12029_ VPWR VGND _00607_ sg13g2_mux2_1
X_19272_ _12024_ \atbs_core_0.uart_0.uart_tx_0.n3349_o\ VPWR VGND _12050_ sg13g2_nor2b_1
X_19273_ \atbs_core_0.memory2uart_0.n2574_o[1]\ _12034_ _12050_ VPWR VGND _12051_ sg13g2_a21oi_1
X_19274_ _12021_ \atbs_core_0.b_data[17]\ VPWR VGND _12052_ sg13g2_nand2_1
X_19275_ _12022_ _12051_ _12052_ VPWR VGND _00608_ sg13g2_o21ai_1
X_19276_ \atbs_core_0.memory2uart_0.n2574_o[12]\ \atbs_core_0.b_data[4]\ _12029_ VPWR VGND _00609_ sg13g2_mux2_1
X_19277_ \atbs_core_0.memory2uart_0.n2574_o[13]\ \atbs_core_0.b_data[5]\ _12029_ VPWR VGND _00610_ sg13g2_mux2_1
X_19278_ \atbs_core_0.memory2uart_0.n2574_o[14]\ \atbs_core_0.b_data[6]\ _12029_ VPWR VGND _00611_ sg13g2_mux2_1
X_19279_ \atbs_core_0.memory2uart_0.n2574_o[15]\ \atbs_core_0.b_data[7]\ _12029_ VPWR VGND _00612_ sg13g2_mux2_1
X_19280_ \atbs_core_0.memory2uart_0.n2574_o[2]\ _12034_ VPWR VGND _12053_ sg13g2_nand2b_1
X_19281_ \atbs_core_0.uart_0.uart_tx_0.n3350_o\ _12025_ _12053_ VPWR VGND _12054_ sg13g2_o21ai_1
X_19282_ _12020_ \atbs_core_0.b_data[18]\ VPWR VGND _12055_ sg13g2_nor2_1
X_19283_ _12055_ VPWR VGND _12056_ sg13g2_buf_1
X_19284_ _12020_ _12054_ _12056_ VPWR VGND _00613_ sg13g2_a21oi_1
X_19285_ \atbs_core_0.memory2uart_0.n2574_o[3]\ _12034_ VPWR VGND _12057_ sg13g2_nand2b_1
X_19286_ \atbs_core_0.uart_0.uart_tx_0.n3351_o\ _12025_ _12057_ VPWR VGND _12058_ sg13g2_o21ai_1
X_19287_ _12020_ _12058_ _12056_ VPWR VGND _00614_ sg13g2_a21oi_1
X_19288_ \atbs_core_0.memory2uart_0.n2574_o[4]\ _12026_ VPWR VGND _12059_ sg13g2_nand2b_1
X_19289_ \atbs_core_0.uart_0.uart_tx_0.n3352_o\ _12025_ _12059_ VPWR VGND _12060_ sg13g2_o21ai_1
X_19290_ _12020_ _12060_ _12056_ VPWR VGND _00615_ sg13g2_a21oi_1
X_19291_ \atbs_core_0.memory2uart_0.n2574_o[5]\ _12026_ VPWR VGND _12061_ sg13g2_nand2b_1
X_19292_ \atbs_core_0.uart_0.uart_tx_0.n3353_o\ _12025_ _12061_ VPWR VGND _12062_ sg13g2_o21ai_1
X_19293_ _12020_ _12062_ _12056_ VPWR VGND _00616_ sg13g2_a21oi_1
X_19294_ \atbs_core_0.memory2uart_0.n2574_o[6]\ _12026_ VPWR VGND _12063_ sg13g2_nand2b_1
X_19295_ \atbs_core_0.uart_0.uart_tx_0.n3354_o\ _12025_ _12063_ VPWR VGND _12064_ sg13g2_o21ai_1
X_19296_ _12020_ _12064_ _12056_ VPWR VGND _00617_ sg13g2_a21oi_1
X_19297_ \atbs_core_0.memory2uart_0.n2574_o[7]\ _12026_ VPWR VGND _12065_ sg13g2_nand2b_1
X_19298_ \atbs_core_0.uart_0.uart_tx_0.n3355_o\ _12025_ _12065_ VPWR VGND _12066_ sg13g2_o21ai_1
X_19299_ _12020_ _12066_ _12056_ VPWR VGND _00618_ sg13g2_a21oi_1
X_19300_ _12024_ \atbs_core_0.memory2uart_0.n2574_o[0]\ VPWR VGND _12067_ sg13g2_nor2b_1
X_19301_ \atbs_core_0.memory2uart_0.n2574_o[8]\ _12034_ _12067_ VPWR VGND _12068_ sg13g2_a21oi_1
X_19302_ _12021_ \atbs_core_0.b_data[8]\ VPWR VGND _12069_ sg13g2_nand2_1
X_19303_ _12022_ _12068_ _12069_ VPWR VGND _00619_ sg13g2_o21ai_1
X_19304_ _12024_ \atbs_core_0.memory2uart_0.n2574_o[1]\ VPWR VGND _12070_ sg13g2_nor2b_1
X_19305_ \atbs_core_0.memory2uart_0.n2574_o[9]\ _12034_ _12070_ VPWR VGND _12071_ sg13g2_a21oi_1
X_19306_ _12021_ \atbs_core_0.b_data[9]\ VPWR VGND _12072_ sg13g2_nand2_1
X_19307_ _12022_ _12071_ _12072_ VPWR VGND _00620_ sg13g2_o21ai_1
X_19308_ _12025_ _12018_ \atbs_core_0.memory2uart_0.counter[0]\ VPWR VGND _00621_ sg13g2_mux2_1
X_19309_ _12017_ \atbs_core_0.memory2uart_0.counter[1]\ VPWR VGND _12073_ sg13g2_nor2b_1
X_19310_ \atbs_core_0.memory2uart_0.counter[0]\ _12025_ _12073_ VPWR VGND _00622_ sg13g2_a21o_1
X_19311_ _08009_ _07681_ \atbs_core_0.detection_en\ VPWR VGND _12074_ sg13g2_o21ai_1
X_19312_ _07992_ _12074_ VPWR VGND _00623_ sg13g2_nand2_1
X_19313_ _07684_ _07905_ VPWR VGND _12075_ sg13g2_nor2_1
X_19314_ \atbs_core_0.clear_dac\ _07709_ VPWR VGND _12076_ sg13g2_nor2_1
X_19315_ _12075_ _12076_ VPWR VGND _00624_ sg13g2_nor2_1
X_19316_ _07541_ _07547_ VPWR VGND _12077_ sg13g2_or2_1
X_19317_ _12077_ VPWR VGND _12078_ sg13g2_buf_1
X_19318_ _12078_ VPWR VGND _12079_ sg13g2_buf_1
X_19319_ _07523_ _07522_ VPWR VGND _12080_ sg13g2_xor2_1
X_19320_ _12080_ _07560_ VPWR VGND _12081_ sg13g2_nand2_1
X_19321_ _07528_ _07558_ VPWR VGND _12082_ sg13g2_nand2_1
X_19322_ _12081_ _12082_ VPWR VGND _12083_ sg13g2_and2_1
X_19323_ _12083_ VPWR VGND _12084_ sg13g2_buf_1
X_19324_ _12084_ VPWR VGND _12085_ sg13g2_buf_1
X_19325_ _12085_ VPWR VGND _12086_ sg13g2_buf_1
X_19326_ _12086_ VPWR VGND _12087_ sg13g2_buf_1
X_19327_ _12087_ VPWR VGND _12088_ sg13g2_buf_1
X_19328_ _07530_ _07550_ VPWR VGND _12089_ sg13g2_xor2_1
X_19329_ _12089_ VPWR VGND _12090_ sg13g2_buf_1
X_19330_ _07533_ _07553_ VPWR VGND _12091_ sg13g2_xnor2_1
X_19331_ _12090_ _12091_ VPWR VGND _12092_ sg13g2_nand2_1
X_19332_ _12092_ VPWR VGND _12093_ sg13g2_buf_1
X_19333_ _12093_ VPWR VGND _12094_ sg13g2_buf_1
X_19334_ _12094_ VPWR VGND _12095_ sg13g2_buf_1
X_19335_ _07909_ _07681_ _07903_ VPWR VGND _12096_ sg13g2_nand3_1
X_19336_ _12096_ VPWR VGND _12097_ sg13g2_buf_1
X_19337_ _12079_ _12088_ _12095_ _12097_ VPWR VGND 
+ _12098_
+ sg13g2_nor4_1
X_19338_ _07903_ _07914_ VPWR VGND _12099_ sg13g2_nand2b_1
X_19339_ _07681_ _12099_ \atbs_core_0.n1389_q\ VPWR VGND _12100_ sg13g2_a21oi_1
X_19340_ _07681_ \atbs_core_0.n1389_q\ _08009_ VPWR VGND _12101_ sg13g2_a21oi_1
X_19341_ _12098_ _12100_ _12101_ VPWR VGND _00625_ sg13g2_nor3_1
X_19342_ _07564_ VPWR VGND _12102_ sg13g2_inv_1
X_19343_ _00056_ _07905_ _07681_ VPWR VGND _12103_ sg13g2_a21oi_1
X_19344_ _12102_ _12103_ \atbs_core_0.enable_read\ VPWR VGND _12104_ sg13g2_o21ai_1
X_19345_ _07564_ _12097_ _12104_ VPWR VGND _00626_ sg13g2_o21ai_1
X_19346_ _07878_ _07879_ VPWR VGND _12105_ sg13g2_nor2_1
X_19347_ _07898_ _12105_ VPWR VGND _12106_ sg13g2_and2_1
X_19348_ _12106_ VPWR VGND _12107_ sg13g2_buf_1
X_19349_ _07877_ _12107_ VPWR VGND _12108_ sg13g2_nand2_1
X_19350_ _07877_ _07886_ VPWR VGND _12109_ sg13g2_nand2_1
X_19351_ _07865_ _07866_ _07856_ _07857_ VPWR VGND 
+ _12110_
+ sg13g2_nor4_1
X_19352_ _07859_ _07860_ VPWR VGND _12111_ sg13g2_nor2b_1
X_19353_ _00060_ _12111_ VPWR VGND _12112_ sg13g2_and2_1
X_19354_ _07855_ _12109_ _12110_ _12112_ VPWR VGND 
+ _12113_
+ sg13g2_nand4_1
X_19355_ _07860_ _07859_ VPWR VGND _12114_ sg13g2_nand2b_1
X_19356_ _12108_ _12113_ _12114_ VPWR VGND _00627_ sg13g2_o21ai_1
X_19357_ _07859_ _07860_ VPWR VGND _12115_ sg13g2_nand2_1
X_19358_ _07872_ _07875_ VPWR VGND _12116_ sg13g2_nor2_1
X_19359_ _07871_ _12116_ VPWR VGND _12117_ sg13g2_nand2_1
X_19360_ _07881_ _07882_ _12105_ _12117_ VPWR VGND 
+ _12118_
+ sg13g2_nor4_1
X_19361_ _12118_ VPWR VGND _12119_ sg13g2_buf_1
X_19362_ _07871_ _12116_ VPWR VGND _12120_ sg13g2_and2_1
X_19363_ _12120_ VPWR VGND _12121_ sg13g2_buf_1
X_19364_ _12107_ _12121_ VPWR VGND _12122_ sg13g2_and2_1
X_19365_ _12122_ VPWR VGND _12123_ sg13g2_buf_1
X_19366_ _12119_ _12123_ VPWR VGND _12124_ sg13g2_nor2_1
X_19367_ _07896_ _07898_ _12121_ VPWR VGND _12125_ sg13g2_and3_1
X_19368_ _12125_ VPWR VGND _12126_ sg13g2_buf_1
X_19369_ _12126_ VPWR VGND _12127_ sg13g2_inv_1
X_19370_ _12127_ _12115_ \atbs_core_0.analog_trigger_0.period_adj_i[3]\ VPWR VGND _12128_ sg13g2_o21ai_1
X_19371_ _12115_ _12124_ _12128_ VPWR VGND _00628_ sg13g2_o21ai_1
X_19372_ _12105_ _12121_ _07884_ VPWR VGND _12129_ sg13g2_nand3b_1
X_19373_ _12129_ VPWR VGND _12130_ sg13g2_buf_1
X_19374_ _12119_ _12123_ VPWR VGND _12131_ sg13g2_or2_1
X_19375_ _12131_ VPWR VGND _12132_ sg13g2_buf_1
X_19376_ _12126_ _12132_ VPWR VGND _12133_ sg13g2_nor2_1
X_19377_ _12115_ _12133_ \atbs_core_0.analog_trigger_0.period_adj_i[4]\ VPWR VGND _12134_ sg13g2_o21ai_1
X_19378_ _12115_ _12130_ _12134_ VPWR VGND _00629_ sg13g2_o21ai_1
X_19379_ _07886_ _12121_ VPWR VGND _12135_ sg13g2_nand2_1
X_19380_ _07884_ _07896_ _12121_ VPWR VGND _12136_ sg13g2_nand3_1
X_19381_ _12136_ VPWR VGND _12137_ sg13g2_buf_1
X_19382_ _12135_ _12137_ VPWR VGND _12138_ sg13g2_nand2_1
X_19383_ _12138_ VPWR VGND _12139_ sg13g2_buf_1
X_19384_ _12115_ _12133_ VPWR VGND _12140_ sg13g2_nor2_1
X_19385_ \atbs_core_0.analog_trigger_0.period_adj_i[5]\ _12139_ _12140_ VPWR VGND _00630_ sg13g2_mux2_1
X_19386_ _07884_ _07896_ _12121_ VPWR VGND _12141_ sg13g2_and3_1
X_19387_ _12141_ VPWR VGND _12142_ sg13g2_buf_1
X_19388_ \atbs_core_0.analog_trigger_0.period_adj_i[6]\ _12142_ _12140_ VPWR VGND _00631_ sg13g2_mux2_1
X_19389_ _07871_ _07872_ _07875_ VPWR VGND _12143_ sg13g2_nor3_1
X_19390_ _12143_ VPWR VGND _12144_ sg13g2_buf_1
X_19391_ _07878_ _07880_ _07898_ _12144_ VPWR VGND 
+ _12145_
+ sg13g2_nand4_1
X_19392_ _07858_ _07861_ VPWR VGND _12146_ sg13g2_nand2_1
X_19393_ _12113_ _12145_ _12146_ VPWR VGND _00632_ sg13g2_o21ai_1
X_19394_ _07858_ _12111_ VPWR VGND _12147_ sg13g2_and2_1
X_19395_ _12147_ VPWR VGND _12148_ sg13g2_buf_1
X_19396_ _12119_ _12148_ _00164_ VPWR VGND _12149_ sg13g2_a21oi_1
X_19397_ _12139_ _12148_ _12149_ VPWR VGND _00633_ sg13g2_a21oi_1
X_19398_ \atbs_core_0.n1394_q[7]\ VPWR VGND _12150_ sg13g2_buf_1
X_19399_ _12150_ VPWR VGND _12151_ sg13g2_inv_1
X_19400_ _12119_ _12148_ _12151_ VPWR VGND _12152_ sg13g2_a21oi_1
X_19401_ _12142_ _12148_ _12152_ VPWR VGND _00634_ sg13g2_a21o_1
X_19402_ _00066_ _07862_ _07867_ VPWR VGND _12153_ sg13g2_and3_1
X_19403_ _12153_ VPWR VGND _12154_ sg13g2_buf_1
X_19404_ _07855_ _12144_ _12154_ VPWR VGND _12155_ sg13g2_nand3_1
X_19405_ _07881_ _07882_ VPWR VGND _12156_ sg13g2_nor2b_1
X_19406_ _07896_ _12156_ VPWR VGND _12157_ sg13g2_nand2_1
X_19407_ _07858_ _07861_ _07857_ VPWR VGND _12158_ sg13g2_o21ai_1
X_19408_ _12155_ _12157_ _12158_ VPWR VGND _00635_ sg13g2_o21ai_1
X_19409_ _07857_ _12112_ VPWR VGND _12159_ sg13g2_and2_1
X_19410_ _12159_ VPWR VGND _12160_ sg13g2_buf_1
X_19411_ _12119_ _12160_ _00165_ VPWR VGND _12161_ sg13g2_a21oi_1
X_19412_ _12139_ _12160_ _12161_ VPWR VGND _00636_ sg13g2_a21oi_1
X_19413_ \atbs_core_0.n1396_q[7]\ VPWR VGND _12162_ sg13g2_buf_1
X_19414_ _12162_ VPWR VGND _12163_ sg13g2_inv_1
X_19415_ _12119_ _12160_ _12163_ VPWR VGND _12164_ sg13g2_a21oi_1
X_19416_ _12142_ _12160_ _12164_ VPWR VGND _00637_ sg13g2_a21o_1
X_19417_ _07862_ _07856_ VPWR VGND _12165_ sg13g2_nand2b_1
X_19418_ _07910_ _12155_ _12165_ VPWR VGND _00638_ sg13g2_o21ai_1
X_19419_ _07856_ _07862_ VPWR VGND _12166_ sg13g2_nand2_1
X_19420_ _12166_ VPWR VGND _12167_ sg13g2_inv_1
X_19421_ _12119_ _12167_ _00166_ VPWR VGND _12168_ sg13g2_a21oi_1
X_19422_ _12139_ _12167_ _12168_ VPWR VGND _00639_ sg13g2_a21oi_1
X_19423_ \atbs_core_0.n1398_q[7]\ VPWR VGND _12169_ sg13g2_buf_1
X_19424_ _12130_ _12166_ _12169_ VPWR VGND _12170_ sg13g2_o21ai_1
X_19425_ _12137_ _12166_ _12170_ VPWR VGND _00640_ sg13g2_o21ai_1
X_19426_ _07895_ _07880_ _07898_ _12144_ VPWR VGND 
+ _12171_
+ sg13g2_nand4_1
X_19427_ _07880_ _07898_ VPWR VGND _12172_ sg13g2_nand2_1
X_19428_ _07880_ _12156_ VPWR VGND _12173_ sg13g2_nand2b_1
X_19429_ _12172_ _12173_ _07895_ VPWR VGND _12174_ sg13g2_a21oi_1
X_19430_ _07880_ _12105_ _07881_ VPWR VGND _12175_ sg13g2_mux2_1
X_19431_ _07882_ _07877_ _12175_ VPWR VGND _12176_ sg13g2_nand3b_1
X_19432_ _07866_ _07864_ VPWR VGND _12177_ sg13g2_nor2b_1
X_19433_ _00107_ _07855_ _12176_ _12177_ VPWR VGND 
+ _12178_
+ sg13g2_nand4_1
X_19434_ _12144_ _12174_ _12178_ VPWR VGND _12179_ sg13g2_a21o_1
X_19435_ _07864_ _07866_ VPWR VGND _12180_ sg13g2_nand2b_1
X_19436_ _12171_ _12179_ _12180_ VPWR VGND _00641_ sg13g2_o21ai_1
X_19437_ _07866_ _07864_ VPWR VGND _12181_ sg13g2_nand2_1
X_19438_ \atbs_core_0.n1400_q[10]\ VPWR VGND _12182_ sg13g2_buf_1
X_19439_ _12135_ _12181_ _12182_ VPWR VGND _12183_ sg13g2_o21ai_1
X_19440_ _12137_ _12181_ _12183_ VPWR VGND _00642_ sg13g2_o21ai_1
X_19441_ _07877_ _07884_ _12105_ VPWR VGND _12184_ sg13g2_nand3_1
X_19442_ _12177_ _07865_ VPWR VGND _12185_ sg13g2_nand2b_1
X_19443_ _12179_ _12184_ _12185_ VPWR VGND _00643_ sg13g2_o21ai_1
X_19444_ _07865_ _12132_ _12177_ VPWR VGND _12186_ sg13g2_nand3_1
X_19445_ _12186_ VPWR VGND _12187_ sg13g2_buf_1
X_19446_ _00167_ _12187_ VPWR VGND _12188_ sg13g2_nand2_1
X_19447_ _12119_ _12187_ _12188_ VPWR VGND _00644_ sg13g2_o21ai_1
X_19448_ _00168_ _12187_ VPWR VGND _12189_ sg13g2_nand2_1
X_19449_ _12139_ _12187_ _12189_ VPWR VGND _00645_ sg13g2_o21ai_1
X_19450_ _00169_ _12187_ VPWR VGND _12190_ sg13g2_nand2_1
X_19451_ _12142_ _12187_ _12190_ VPWR VGND _00646_ sg13g2_o21ai_1
X_19452_ _07852_ VPWR VGND _12191_ sg13g2_inv_1
X_19453_ _07895_ _07880_ _07898_ VPWR VGND _12192_ sg13g2_nand3_1
X_19454_ _12192_ VPWR VGND _12193_ sg13g2_buf_1
X_19455_ _07851_ VPWR VGND _12194_ sg13g2_inv_1
X_19456_ _12194_ _00064_ _07850_ _07886_ VPWR VGND 
+ _12195_
+ sg13g2_and4_1
X_19457_ _12144_ _12154_ _12193_ _12195_ VPWR VGND 
+ _12196_
+ sg13g2_nand4_1
X_19458_ _12191_ _12154_ _12196_ VPWR VGND _00647_ sg13g2_o21ai_1
X_19459_ _07852_ _12154_ VPWR VGND _12197_ sg13g2_nand2_1
X_19460_ _12197_ _12132_ VPWR VGND _12198_ sg13g2_nand2b_1
X_19461_ _12198_ VPWR VGND _12199_ sg13g2_buf_1
X_19462_ _00170_ _12199_ VPWR VGND _12200_ sg13g2_nand2_1
X_19463_ _12135_ _12199_ _12200_ VPWR VGND _00648_ sg13g2_o21ai_1
X_19464_ _12130_ _12197_ VPWR VGND _12201_ sg13g2_nor2_1
X_19465_ _00171_ _12199_ _12201_ VPWR VGND _00649_ sg13g2_a21o_1
X_19466_ _07910_ _12121_ VPWR VGND _12202_ sg13g2_nand2b_1
X_19467_ _07585_ _12199_ VPWR VGND _12203_ sg13g2_nand2_1
X_19468_ _12197_ _12202_ _12203_ VPWR VGND _00650_ sg13g2_o21ai_1
X_19469_ _07590_ _12199_ VPWR VGND _12204_ sg13g2_nand2_1
X_19470_ _12135_ _12199_ _12204_ VPWR VGND _00651_ sg13g2_o21ai_1
X_19471_ _07580_ VPWR VGND _12205_ sg13g2_inv_1
X_19472_ _12124_ _12197_ VPWR VGND _12206_ sg13g2_nor2_1
X_19473_ _12142_ _12206_ VPWR VGND _12207_ sg13g2_nand2_1
X_19474_ _12205_ _12206_ _12207_ VPWR VGND _00652_ sg13g2_o21ai_1
X_19475_ _07878_ _07884_ _12121_ VPWR VGND _12208_ sg13g2_nand3_1
X_19476_ _00172_ _12199_ VPWR VGND _12209_ sg13g2_nand2_1
X_19477_ _12199_ _12208_ _12209_ VPWR VGND _00653_ sg13g2_o21ai_1
X_19478_ _07569_ _12199_ _12201_ VPWR VGND _00654_ sg13g2_a21o_1
X_19479_ _07894_ _12193_ VPWR VGND _12210_ sg13g2_nor2_1
X_19480_ _07852_ _07900_ VPWR VGND _12211_ sg13g2_nor2_1
X_19481_ _07851_ _12210_ _12211_ VPWR VGND _00655_ sg13g2_mux2_1
X_19482_ _07851_ _12132_ _12211_ VPWR VGND _12212_ sg13g2_nand3_1
X_19483_ _12212_ VPWR VGND _12213_ sg13g2_buf_1
X_19484_ _11423_ _12213_ VPWR VGND _12214_ sg13g2_nand2_1
X_19485_ _12137_ _12213_ _12214_ VPWR VGND _00656_ sg13g2_o21ai_1
X_19486_ _07886_ _12121_ VPWR VGND _12215_ sg13g2_and2_1
X_19487_ _00173_ _12213_ VPWR VGND _12216_ sg13g2_nand2_1
X_19488_ _12215_ _12213_ _12216_ VPWR VGND _00657_ sg13g2_o21ai_1
X_19489_ _11395_ _12213_ VPWR VGND _12217_ sg13g2_nand2_1
X_19490_ _12202_ _12213_ _12217_ VPWR VGND _00658_ sg13g2_o21ai_1
X_19491_ _11386_ _12213_ VPWR VGND _12218_ sg13g2_nand2_1
X_19492_ _12119_ _12213_ _12218_ VPWR VGND _00659_ sg13g2_o21ai_1
X_19493_ _00108_ _07877_ VPWR VGND _12219_ sg13g2_nand2_1
X_19494_ _07895_ _07849_ _12172_ _12219_ VPWR VGND 
+ _12220_
+ sg13g2_nor4_1
X_19495_ _07853_ _12154_ VPWR VGND _12221_ sg13g2_nand2_1
X_19496_ _12220_ _07849_ _12221_ VPWR VGND _00660_ sg13g2_mux2_1
X_19497_ _12126_ _12119_ VPWR VGND _12222_ sg13g2_nor2_1
X_19498_ _12117_ _12193_ _12133_ VPWR VGND _12223_ sg13g2_o21ai_1
X_19499_ _07849_ _07853_ _12154_ _12223_ VPWR VGND 
+ _12224_
+ sg13g2_and4_1
X_19500_ _12224_ VPWR VGND _12225_ sg13g2_buf_1
X_19501_ _12225_ VPWR VGND _12226_ sg13g2_buf_1
X_19502_ _00174_ _12222_ _12226_ VPWR VGND _00661_ sg13g2_mux2_1
X_19503_ _00175_ _12126_ _12226_ VPWR VGND _00662_ sg13g2_mux2_1
X_19504_ _00176_ VPWR VGND _12227_ sg13g2_inv_1
X_19505_ _12133_ _12225_ VPWR VGND _12228_ sg13g2_nand2_1
X_19506_ _12227_ _12226_ _12228_ VPWR VGND _00663_ sg13g2_o21ai_1
X_19507_ _00177_ VPWR VGND _12229_ sg13g2_inv_1
X_19508_ _12142_ _12225_ VPWR VGND _12230_ sg13g2_nand2_1
X_19509_ _12229_ _12226_ _12230_ VPWR VGND _00664_ sg13g2_o21ai_1
X_19510_ _00178_ _12139_ _12225_ VPWR VGND _00665_ sg13g2_mux2_1
X_19511_ _12130_ _12225_ VPWR VGND _12231_ sg13g2_nand2_1
X_19512_ _08696_ _12226_ _12231_ VPWR VGND _00666_ sg13g2_o21ai_1
X_19513_ _12124_ _12225_ VPWR VGND _12232_ sg13g2_nand2_1
X_19514_ _08716_ _12226_ _12232_ VPWR VGND _00667_ sg13g2_o21ai_1
X_19515_ _08712_ _12226_ _12228_ VPWR VGND _00668_ sg13g2_o21ai_1
X_19516_ _08516_ _12226_ _12230_ VPWR VGND _00669_ sg13g2_o21ai_1
X_19517_ _12215_ _12225_ VPWR VGND _12233_ sg13g2_nand2_1
X_19518_ _09361_ _12226_ _12233_ VPWR VGND _00670_ sg13g2_o21ai_1
X_19519_ _00179_ _12208_ _12225_ VPWR VGND _00671_ sg13g2_mux2_1
X_19520_ _12123_ _12139_ _12225_ VPWR VGND _12234_ sg13g2_o21ai_1
X_19521_ _08625_ _12226_ _12234_ VPWR VGND _00672_ sg13g2_o21ai_1
X_19522_ _00108_ _12107_ _12144_ _12193_ VPWR VGND 
+ _12235_
+ sg13g2_and4_1
X_19523_ _07849_ _07851_ _07852_ _07900_ VPWR VGND 
+ _12236_
+ sg13g2_nor4_1
X_19524_ \atbs_core_0.atbs_max_delta_steps_uart\ _12235_ _12236_ VPWR VGND _00673_ sg13g2_mux2_1
X_19525_ _07849_ \atbs_core_0.atbs_max_delta_steps_uart\ VPWR VGND _12237_ sg13g2_nor2b_1
X_19526_ _07853_ _07868_ _12132_ _12237_ VPWR VGND 
+ _12238_
+ sg13g2_nand4_1
X_19527_ _12238_ VPWR VGND _12239_ sg13g2_buf_1
X_19528_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[1]\ _12239_ VPWR VGND _12240_ sg13g2_nand2_1
X_19529_ _12137_ _12239_ _12240_ VPWR VGND _00674_ sg13g2_o21ai_1
X_19530_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _12239_ VPWR VGND _12241_ sg13g2_nand2_1
X_19531_ _12135_ _12239_ _12241_ VPWR VGND _00675_ sg13g2_o21ai_1
X_19532_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _12239_ VPWR VGND _12242_ sg13g2_nand2_1
X_19533_ _12202_ _12239_ _12242_ VPWR VGND _00676_ sg13g2_o21ai_1
X_19534_ _00180_ _12239_ VPWR VGND _12243_ sg13g2_nand2_1
X_19535_ _12130_ _12239_ _12243_ VPWR VGND _00677_ sg13g2_o21ai_1
X_19536_ _07909_ _07903_ _07680_ _07684_ VPWR VGND 
+ _12244_
+ sg13g2_nor4_1
X_19537_ _07680_ _07902_ VPWR VGND _12245_ sg13g2_and2_1
X_19538_ _07906_ _12245_ idle_led_o VPWR VGND _12246_ sg13g2_a21oi_1
X_19539_ _12244_ _12246_ VPWR VGND _00678_ sg13g2_nor2_1
X_19540_ overflow_led_o _12098_ VPWR VGND _12247_ sg13g2_nor2_1
X_19541_ _12075_ _12247_ VPWR VGND _00679_ sg13g2_nor2_1
X_19542_ _12078_ _12084_ _12093_ VPWR VGND _12248_ sg13g2_nor3_1
X_19543_ _12248_ _12097_ VPWR VGND _12249_ sg13g2_nor2_1
X_19544_ underflow_led_o _07564_ _12249_ VPWR VGND _12250_ sg13g2_mux2_1
X_19545_ _12075_ _12250_ VPWR VGND _00680_ sg13g2_nor2b_1
X_19546_ \atbs_core_0.uart_0.uart_rx_0.n3486_o\ \atbs_core_0.uart_0.uart_rx_0.n3484_o\ VPWR VGND _12251_ sg13g2_nor2_1
X_19547_ _07871_ _07872_ _07870_ _12251_ VPWR VGND 
+ _12252_
+ sg13g2_nand4_1
X_19548_ _12252_ VPWR VGND _12253_ sg13g2_buf_1
X_19549_ _07880_ _12253_ VPWR VGND _12254_ sg13g2_nor2_1
X_19550_ _07884_ _12254_ VPWR VGND _12255_ sg13g2_nand2_1
X_19551_ _00181_ _12255_ VPWR VGND _12256_ sg13g2_nand2_1
X_19552_ _07878_ _12255_ _12256_ VPWR VGND _00681_ sg13g2_o21ai_1
X_19553_ _07885_ _12253_ VPWR VGND _12257_ sg13g2_nor2_1
X_19554_ \atbs_core_0.adaptive_mode_uart\ _07878_ _12257_ VPWR VGND _00682_ sg13g2_mux2_1
X_19555_ _07898_ _12254_ VPWR VGND _12258_ sg13g2_nand2_1
X_19556_ _00182_ _12258_ VPWR VGND _12259_ sg13g2_nand2_1
X_19557_ _07878_ _12258_ _12259_ VPWR VGND _00683_ sg13g2_o21ai_1
X_19558_ _12172_ _12253_ VPWR VGND _12260_ sg13g2_nor2_1
X_19559_ _00183_ _07895_ _12260_ VPWR VGND _00684_ sg13g2_mux2_1
X_19560_ _12156_ _12254_ VPWR VGND _12261_ sg13g2_nand2_1
X_19561_ _00184_ _12261_ VPWR VGND _12262_ sg13g2_nand2_1
X_19562_ _07878_ _12261_ _12262_ VPWR VGND _00685_ sg13g2_o21ai_1
X_19563_ \atbs_core_0.sc_noc_generator_0.counter_value[0]\ VPWR VGND _12263_ sg13g2_buf_1
X_19564_ _12263_ _07680_ VPWR VGND _00686_ sg13g2_xnor2_1
X_19565_ \atbs_core_0.sc_noc_generator_0.counter_value[1]\ VPWR VGND _12264_ sg13g2_buf_1
X_19566_ _12263_ _07658_ VPWR VGND _12265_ sg13g2_nand2_1
X_19567_ _12264_ _12265_ VPWR VGND _00687_ sg13g2_xnor2_1
X_19568_ \atbs_core_0.sc_noc_generator_0.counter_value[2]\ VPWR VGND _12266_ sg13g2_buf_1
X_19569_ _12264_ _12263_ _07657_ VPWR VGND _12267_ sg13g2_nand3_1
X_19570_ _12266_ _12267_ VPWR VGND _00688_ sg13g2_xnor2_1
X_19571_ _12264_ _12263_ _12266_ _07658_ VPWR VGND 
+ _12268_
+ sg13g2_nand4_1
X_19572_ \atbs_core_0.sc_noc_generator_0.counter_value[3]\ _12268_ VPWR VGND _00689_ sg13g2_xnor2_1
X_19573_ _12266_ \atbs_core_0.sc_noc_generator_0.counter_value[3]\ VPWR VGND _12269_ sg13g2_and2_1
X_19574_ _12267_ _12269_ VPWR VGND _12270_ sg13g2_nand2b_1
X_19575_ \atbs_core_0.sc_noc_generator_0.counter_value[4]\ _12270_ VPWR VGND _00690_ sg13g2_xnor2_1
X_19576_ \atbs_core_0.sc_noc_generator_0.counter_value[5]\ VPWR VGND _12271_ sg13g2_buf_1
X_19577_ _12264_ \atbs_core_0.sc_noc_generator_0.counter_value[4]\ _12269_ VPWR VGND _12272_ sg13g2_and3_1
X_19578_ _12263_ _12272_ VPWR VGND _12273_ sg13g2_and2_1
X_19579_ _12273_ VPWR VGND _12274_ sg13g2_buf_1
X_19580_ _07658_ _12274_ VPWR VGND _12275_ sg13g2_nand2_1
X_19581_ _12271_ _12275_ VPWR VGND _00691_ sg13g2_xnor2_1
X_19582_ _00034_ VPWR VGND _12276_ sg13g2_buf_1
X_19583_ _12150_ \atbs_core_0.sc_noc_generator_0.counter_value[7]\ VPWR VGND _12277_ sg13g2_xnor2_1
X_19584_ \atbs_core_0.sc_noc_generator_0.counter_value[6]\ VPWR VGND _12278_ sg13g2_buf_1
X_19585_ \atbs_core_0.n1394_q[6]\ VPWR VGND _12279_ sg13g2_buf_1
X_19586_ _12278_ _12279_ VPWR VGND _12280_ sg13g2_xnor2_1
X_19587_ _12277_ _12280_ VPWR VGND _12281_ sg13g2_nand2_1
X_19588_ _12276_ _12281_ VPWR VGND _12282_ sg13g2_nand2_1
X_19589_ _12271_ _12274_ VPWR VGND _12283_ sg13g2_nand2_1
X_19590_ _12282_ _12276_ _12283_ VPWR VGND _12284_ sg13g2_mux2_1
X_19591_ _12278_ _07844_ VPWR VGND _12285_ sg13g2_nor2_1
X_19592_ bio_amp_en_o _12284_ _12285_ VPWR VGND _00692_ sg13g2_a21oi_1
X_19593_ _00035_ VPWR VGND _12286_ sg13g2_buf_1
X_19594_ _12286_ VPWR VGND _12287_ sg13g2_inv_1
X_19595_ _12271_ _12278_ _12286_ _12274_ VPWR VGND 
+ _12288_
+ sg13g2_nand4_1
X_19596_ _12278_ _12286_ _12288_ VPWR VGND _12289_ sg13g2_o21ai_1
X_19597_ _12287_ _12283_ _12281_ _12289_ VPWR VGND 
+ _12290_
+ sg13g2_a22oi_1
X_19598_ \atbs_core_0.sc_noc_generator_0.counter_value[7]\ _07844_ VPWR VGND _12291_ sg13g2_nor2_1
X_19599_ bio_amp_en_o _12290_ _12291_ VPWR VGND _00693_ sg13g2_a21oi_1
X_19600_ \atbs_core_0.sc_noc_generator_1.counter_value[0]\ VPWR VGND _12292_ sg13g2_buf_1
X_19601_ _12292_ _07680_ VPWR VGND _00694_ sg13g2_xnor2_1
X_19602_ \atbs_core_0.sc_noc_generator_1.counter_value[1]\ VPWR VGND _12293_ sg13g2_buf_1
X_19603_ _12292_ _07658_ VPWR VGND _12294_ sg13g2_nand2_1
X_19604_ _12293_ _12294_ VPWR VGND _00695_ sg13g2_xnor2_1
X_19605_ \atbs_core_0.sc_noc_generator_1.counter_value[2]\ VPWR VGND _12295_ sg13g2_buf_1
X_19606_ _12293_ _12292_ _07657_ VPWR VGND _12296_ sg13g2_nand3_1
X_19607_ _12295_ _12296_ VPWR VGND _00696_ sg13g2_xnor2_1
X_19608_ _12293_ _12292_ _12295_ _07658_ VPWR VGND 
+ _12297_
+ sg13g2_nand4_1
X_19609_ \atbs_core_0.sc_noc_generator_1.counter_value[3]\ _12297_ VPWR VGND _00697_ sg13g2_xnor2_1
X_19610_ \atbs_core_0.sc_noc_generator_1.counter_value[3]\ _12295_ VPWR VGND _12298_ sg13g2_and2_1
X_19611_ _12296_ _12298_ VPWR VGND _12299_ sg13g2_nand2b_1
X_19612_ \atbs_core_0.sc_noc_generator_1.counter_value[4]\ _12299_ VPWR VGND _00698_ sg13g2_xnor2_1
X_19613_ \atbs_core_0.sc_noc_generator_1.counter_value[5]\ VPWR VGND _12300_ sg13g2_buf_1
X_19614_ _12293_ \atbs_core_0.sc_noc_generator_1.counter_value[4]\ _12298_ VPWR VGND _12301_ sg13g2_and3_1
X_19615_ _12292_ _12301_ VPWR VGND _12302_ sg13g2_and2_1
X_19616_ _12302_ VPWR VGND _12303_ sg13g2_buf_1
X_19617_ _07658_ _12303_ VPWR VGND _12304_ sg13g2_nand2_1
X_19618_ _12300_ _12304_ VPWR VGND _00699_ sg13g2_xnor2_1
X_19619_ _00032_ VPWR VGND _12305_ sg13g2_buf_1
X_19620_ _12162_ \atbs_core_0.sc_noc_generator_1.counter_value[7]\ VPWR VGND _12306_ sg13g2_xnor2_1
X_19621_ \atbs_core_0.sc_noc_generator_1.counter_value[6]\ VPWR VGND _12307_ sg13g2_buf_1
X_19622_ \atbs_core_0.n1396_q[6]\ VPWR VGND _12308_ sg13g2_buf_1
X_19623_ _12307_ _12308_ VPWR VGND _12309_ sg13g2_xnor2_1
X_19624_ _12306_ _12309_ VPWR VGND _12310_ sg13g2_nand2_1
X_19625_ _12305_ _12310_ VPWR VGND _12311_ sg13g2_nand2_1
X_19626_ _12300_ _12303_ VPWR VGND _12312_ sg13g2_nand2_1
X_19627_ _12311_ _12305_ _12312_ VPWR VGND _12313_ sg13g2_mux2_1
X_19628_ _12307_ _07844_ VPWR VGND _12314_ sg13g2_nor2_1
X_19629_ bio_amp_en_o _12313_ _12314_ VPWR VGND _00700_ sg13g2_a21oi_1
X_19630_ _00033_ VPWR VGND _12315_ sg13g2_buf_1
X_19631_ _12315_ VPWR VGND _12316_ sg13g2_inv_1
X_19632_ _12300_ _12307_ _12315_ _12303_ VPWR VGND 
+ _12317_
+ sg13g2_nand4_1
X_19633_ _12307_ _12315_ _12317_ VPWR VGND _12318_ sg13g2_o21ai_1
X_19634_ _12316_ _12312_ _12310_ _12318_ VPWR VGND 
+ _12319_
+ sg13g2_a22oi_1
X_19635_ \atbs_core_0.sc_noc_generator_1.counter_value[7]\ _07844_ VPWR VGND _12320_ sg13g2_nor2_1
X_19636_ bio_amp_en_o _12319_ _12320_ VPWR VGND _00701_ sg13g2_a21oi_1
X_19637_ \atbs_core_0.sc_noc_generator_2.counter_value[0]\ VPWR VGND _12321_ sg13g2_buf_1
X_19638_ _12321_ _07680_ VPWR VGND _00702_ sg13g2_xnor2_1
X_19639_ \atbs_core_0.sc_noc_generator_2.counter_value[1]\ VPWR VGND _12322_ sg13g2_buf_1
X_19640_ _12321_ _07658_ VPWR VGND _12323_ sg13g2_nand2_1
X_19641_ _12322_ _12323_ VPWR VGND _00703_ sg13g2_xnor2_1
X_19642_ \atbs_core_0.sc_noc_generator_2.counter_value[2]\ VPWR VGND _12324_ sg13g2_buf_1
X_19643_ _12322_ _12321_ _07657_ VPWR VGND _12325_ sg13g2_nand3_1
X_19644_ _12324_ _12325_ VPWR VGND _00704_ sg13g2_xnor2_1
X_19645_ _12322_ _12321_ _12324_ _07657_ VPWR VGND 
+ _12326_
+ sg13g2_nand4_1
X_19646_ \atbs_core_0.sc_noc_generator_2.counter_value[3]\ _12326_ VPWR VGND _00705_ sg13g2_xnor2_1
X_19647_ \atbs_core_0.sc_noc_generator_2.counter_value[3]\ _12324_ VPWR VGND _12327_ sg13g2_and2_1
X_19648_ _12325_ _12327_ VPWR VGND _12328_ sg13g2_nand2b_1
X_19649_ \atbs_core_0.sc_noc_generator_2.counter_value[4]\ _12328_ VPWR VGND _00706_ sg13g2_xnor2_1
X_19650_ \atbs_core_0.sc_noc_generator_2.counter_value[5]\ VPWR VGND _12329_ sg13g2_buf_1
X_19651_ _12322_ _12321_ \atbs_core_0.sc_noc_generator_2.counter_value[4]\ _12327_ VPWR VGND 
+ _12330_
+ sg13g2_and4_1
X_19652_ _12330_ VPWR VGND _12331_ sg13g2_buf_1
X_19653_ _07658_ _12331_ VPWR VGND _12332_ sg13g2_nand2_1
X_19654_ _12329_ _12332_ VPWR VGND _00707_ sg13g2_xnor2_1
X_19655_ \atbs_core_0.sc_noc_generator_2.counter_value[6]\ VPWR VGND _12333_ sg13g2_buf_1
X_19656_ _00030_ VPWR VGND _12334_ sg13g2_buf_1
X_19657_ _12329_ _12331_ VPWR VGND _12335_ sg13g2_and2_1
X_19658_ _12335_ VPWR VGND _12336_ sg13g2_buf_1
X_19659_ _12169_ \atbs_core_0.sc_noc_generator_2.counter_value[7]\ VPWR VGND _12337_ sg13g2_nor2b_1
X_19660_ _12169_ VPWR VGND _12338_ sg13g2_inv_1
X_19661_ _12338_ \atbs_core_0.sc_noc_generator_2.counter_value[7]\ VPWR VGND _12339_ sg13g2_nor2_1
X_19662_ \atbs_core_0.n1398_q[6]\ VPWR VGND _12340_ sg13g2_buf_1
X_19663_ _12333_ _12340_ VPWR VGND _12341_ sg13g2_xor2_1
X_19664_ _12337_ _12339_ _12341_ VPWR VGND _12342_ sg13g2_or3_1
X_19665_ _12334_ _12336_ _12342_ VPWR VGND _12343_ sg13g2_nand3_1
X_19666_ _12334_ _12336_ _12343_ VPWR VGND _12344_ sg13g2_o21ai_1
X_19667_ _12333_ _12344_ _07844_ VPWR VGND _00708_ sg13g2_mux2_1
X_19668_ _00031_ VPWR VGND _12345_ sg13g2_buf_1
X_19669_ _12345_ VPWR VGND _12346_ sg13g2_inv_1
X_19670_ _12329_ _12331_ VPWR VGND _12347_ sg13g2_nand2_1
X_19671_ _12333_ _12345_ _12336_ VPWR VGND _12348_ sg13g2_nand3_1
X_19672_ _12333_ _12345_ _12348_ VPWR VGND _12349_ sg13g2_o21ai_1
X_19673_ _12346_ _12347_ _12342_ _12349_ VPWR VGND 
+ _12350_
+ sg13g2_a22oi_1
X_19674_ \atbs_core_0.sc_noc_generator_2.counter_value[7]\ _07844_ VPWR VGND _12351_ sg13g2_nor2_1
X_19675_ bio_amp_en_o _12350_ _12351_ VPWR VGND _00709_ sg13g2_a21oi_1
X_19676_ \atbs_core_0.sc_noc_generator_3.counter_value[0]\ VPWR VGND _12352_ sg13g2_buf_1
X_19677_ _12352_ _07680_ VPWR VGND _00710_ sg13g2_xnor2_1
X_19678_ \atbs_core_0.sc_noc_generator_3.counter_value[9]\ VPWR VGND _12353_ sg13g2_buf_1
X_19679_ \atbs_core_0.sc_noc_generator_3.counter_value[8]\ VPWR VGND _12354_ sg13g2_buf_1
X_19680_ \atbs_core_0.sc_noc_generator_3.counter_value[3]\ \atbs_core_0.sc_noc_generator_3.counter_value[5]\ \atbs_core_0.sc_noc_generator_3.counter_value[4]\ VPWR VGND _12355_ sg13g2_nand3_1
X_19681_ \atbs_core_0.sc_noc_generator_3.counter_value[1]\ VPWR VGND _12356_ sg13g2_buf_1
X_19682_ \atbs_core_0.sc_noc_generator_3.counter_value[2]\ VPWR VGND _12357_ sg13g2_buf_1
X_19683_ _12356_ _12357_ \atbs_core_0.sc_noc_generator_3.counter_value[7]\ \atbs_core_0.sc_noc_generator_3.counter_value[6]\ VPWR VGND 
+ _12358_
+ sg13g2_nand4_1
X_19684_ _12355_ _12358_ VPWR VGND _12359_ sg13g2_nor2_1
X_19685_ _12352_ _12354_ _12359_ VPWR VGND _12360_ sg13g2_and3_1
X_19686_ _12360_ VPWR VGND _12361_ sg13g2_buf_1
X_19687_ \atbs_core_0.sc_noc_generator_3.counter_value[10]\ VPWR VGND _12362_ sg13g2_buf_1
X_19688_ _12362_ VPWR VGND _12363_ sg13g2_inv_1
X_19689_ _12182_ _12363_ _07657_ VPWR VGND _12364_ sg13g2_nand3_1
X_19690_ _12182_ _12363_ _12364_ VPWR VGND _12365_ sg13g2_o21ai_1
X_19691_ _12353_ _00029_ _12361_ _12365_ VPWR VGND 
+ _12366_
+ sg13g2_nand4_1
X_19692_ _12353_ _12361_ VPWR VGND _12367_ sg13g2_nand2_1
X_19693_ _00029_ _07680_ VPWR VGND _12368_ sg13g2_nor2_1
X_19694_ _12362_ _07680_ _12367_ _12368_ VPWR VGND 
+ _12369_
+ sg13g2_a22oi_1
X_19695_ _12366_ _12369_ VPWR VGND _00711_ sg13g2_nand2_1
X_19696_ _12352_ _07657_ VPWR VGND _12370_ sg13g2_and2_1
X_19697_ _12370_ VPWR VGND _12371_ sg13g2_buf_1
X_19698_ _12356_ _12371_ VPWR VGND _00712_ sg13g2_xor2_1
X_19699_ _12356_ _12371_ VPWR VGND _12372_ sg13g2_nand2_1
X_19700_ _12357_ _12372_ VPWR VGND _00713_ sg13g2_xnor2_1
X_19701_ _12356_ _12357_ _12371_ VPWR VGND _12373_ sg13g2_nand3_1
X_19702_ \atbs_core_0.sc_noc_generator_3.counter_value[3]\ _12373_ VPWR VGND _00714_ sg13g2_xnor2_1
X_19703_ _12356_ \atbs_core_0.sc_noc_generator_3.counter_value[3]\ _12357_ _12371_ VPWR VGND 
+ _12374_
+ sg13g2_nand4_1
X_19704_ \atbs_core_0.sc_noc_generator_3.counter_value[4]\ _12374_ VPWR VGND _00715_ sg13g2_xnor2_1
X_19705_ \atbs_core_0.sc_noc_generator_3.counter_value[4]\ VPWR VGND _12375_ sg13g2_inv_1
X_19706_ _12375_ _12374_ VPWR VGND _12376_ sg13g2_or2_1
X_19707_ \atbs_core_0.sc_noc_generator_3.counter_value[5]\ _12376_ VPWR VGND _00716_ sg13g2_xnor2_1
X_19708_ _12355_ _12373_ VPWR VGND _12377_ sg13g2_nor2_1
X_19709_ \atbs_core_0.sc_noc_generator_3.counter_value[6]\ _12377_ VPWR VGND _00717_ sg13g2_xor2_1
X_19710_ \atbs_core_0.sc_noc_generator_3.counter_value[6]\ _12377_ VPWR VGND _12378_ sg13g2_nand2_1
X_19711_ \atbs_core_0.sc_noc_generator_3.counter_value[7]\ _12378_ VPWR VGND _00718_ sg13g2_xnor2_1
X_19712_ _12371_ _12359_ VPWR VGND _12379_ sg13g2_nand2_1
X_19713_ _12354_ _12379_ VPWR VGND _00719_ sg13g2_xnor2_1
X_19714_ _12353_ VPWR VGND _12380_ sg13g2_inv_1
X_19715_ _12182_ _12362_ VPWR VGND _12381_ sg13g2_xor2_1
X_19716_ _12380_ _12381_ _00028_ VPWR VGND _12382_ sg13g2_o21ai_1
X_19717_ _00028_ _12382_ _12361_ VPWR VGND _12383_ sg13g2_mux2_1
X_19718_ _12353_ _07844_ VPWR VGND _12384_ sg13g2_nor2_1
X_19719_ bio_amp_en_o _12383_ _12384_ VPWR VGND _00720_ sg13g2_a21oi_1
X_19720_ _07928_ VPWR VGND _12385_ sg13g2_inv_1
X_19721_ _07807_ _12385_ _07716_ VPWR VGND _12386_ sg13g2_a21oi_1
X_19722_ \atbs_core_0.spike_detector_0.is_changing\ _07566_ _11321_ _12386_ VPWR VGND 
+ _00721_
+ sg13g2_a22oi_1
X_19723_ \atbs_core_0.dac_control_0.dac_change_in_progress\ VPWR VGND _12387_ sg13g2_inv_1
X_19724_ _12387_ _11608_ \atbs_core_0.spike_detector_0.n1595_q\ VPWR VGND _12388_ sg13g2_o21ai_1
X_19725_ _07803_ _12388_ VPWR VGND _00722_ sg13g2_nand2_1
X_19726_ _07807_ _08262_ _07802_ VPWR VGND _12389_ sg13g2_a21oi_1
X_19727_ \atbs_core_0.dac_control_1.dac_change_in_progress\ VPWR VGND _12390_ sg13g2_inv_1
X_19728_ _12390_ _11832_ \atbs_core_0.spike_detector_0.lower_is_changing\ VPWR VGND _12391_ sg13g2_o21ai_1
X_19729_ _12389_ _12391_ VPWR VGND _00723_ sg13g2_nand2_1
X_19730_ \atbs_core_0.spike_encoder_0.delayed_spike_strb\ _07921_ _08757_ VPWR VGND _12392_ sg13g2_nor3_1
X_19731_ _12392_ VPWR VGND _12393_ sg13g2_buf_1
X_19732_ _12393_ VPWR VGND \atbs_core_0.spike_encoder_0.n2265_o\ sg13g2_inv_1
X_19733_ _12393_ VPWR VGND _12394_ sg13g2_buf_1
X_19734_ _07921_ _08894_ VPWR VGND _12395_ sg13g2_nand2b_1
X_19735_ \atbs_core_0.encoded_spike[0]\ _12394_ VPWR VGND _12396_ sg13g2_nand2_1
X_19736_ _12394_ _12395_ _12396_ VPWR VGND _00724_ sg13g2_o21ai_1
X_19737_ \atbs_core_0.spike_encoder_0.delayed_spike\ spike_o VPWR VGND _12397_ sg13g2_nor2_1
X_19738_ _12397_ VPWR VGND _12398_ sg13g2_buf_1
X_19739_ _12398_ VPWR VGND _12399_ sg13g2_buf_1
X_19740_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[7]\ VPWR VGND _12400_ sg13g2_buf_1
X_19741_ _08894_ _08892_ _08885_ _08888_ VPWR VGND 
+ _12401_
+ sg13g2_nor4_1
X_19742_ _08884_ _12401_ VPWR VGND _12402_ sg13g2_nand2_1
X_19743_ _08879_ _08557_ _12400_ _12402_ VPWR VGND 
+ _12403_
+ sg13g2_nor4_1
X_19744_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[9]\ VPWR VGND _12404_ sg13g2_buf_1
X_19745_ _10586_ _12404_ VPWR VGND _12405_ sg13g2_nor2_1
X_19746_ _12403_ _12405_ VPWR VGND _12406_ sg13g2_nand2_1
X_19747_ _08860_ _12406_ VPWR VGND _12407_ sg13g2_xnor2_1
X_19748_ _00074_ _12398_ VPWR VGND _12408_ sg13g2_nor2_1
X_19749_ _12399_ _12407_ _12408_ VPWR VGND _12409_ sg13g2_a21oi_1
X_19750_ _07929_ \atbs_core_0.spike_encoder_0.n2265_o\ VPWR VGND _12410_ sg13g2_nand2_1
X_19751_ _12410_ VPWR VGND _12411_ sg13g2_buf_1
X_19752_ _12411_ VPWR VGND _12412_ sg13g2_buf_1
X_19753_ \atbs_core_0.encoded_spike[10]\ _12394_ VPWR VGND _12413_ sg13g2_nand2_1
X_19754_ _12409_ _12412_ _12413_ VPWR VGND _00725_ sg13g2_o21ai_1
X_19755_ _12398_ VPWR VGND _12414_ sg13g2_buf_1
X_19756_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[11]\ VPWR VGND _12415_ sg13g2_buf_1
X_19757_ _12400_ VPWR VGND _12416_ sg13g2_inv_1
X_19758_ _08892_ _00022_ VPWR VGND _12417_ sg13g2_nand2b_1
X_19759_ _12417_ _08889_ _08487_ VPWR VGND _12418_ sg13g2_nand3b_1
X_19760_ _12418_ VPWR VGND _12419_ sg13g2_buf_1
X_19761_ _08879_ _08883_ _08557_ _12419_ VPWR VGND 
+ _12420_
+ sg13g2_nor4_1
X_19762_ _12416_ _12420_ VPWR VGND _12421_ sg13g2_nand2_1
X_19763_ _09048_ _10586_ _12404_ _12421_ VPWR VGND 
+ _12422_
+ sg13g2_nor4_1
X_19764_ _12415_ _12422_ VPWR VGND _12423_ sg13g2_xnor2_1
X_19765_ _12398_ VPWR VGND _12424_ sg13g2_buf_1
X_19766_ _08930_ _12424_ VPWR VGND _12425_ sg13g2_nor2_1
X_19767_ _12414_ _12423_ _12425_ VPWR VGND _12426_ sg13g2_a21oi_1
X_19768_ \atbs_core_0.encoded_spike[11]\ _12394_ VPWR VGND _12427_ sg13g2_nand2_1
X_19769_ _12412_ _12426_ _12427_ VPWR VGND _00726_ sg13g2_o21ai_1
X_19770_ _09048_ _10586_ _12404_ _12415_ VPWR VGND 
+ _12428_
+ sg13g2_nor4_1
X_19771_ _12403_ _12428_ VPWR VGND _12429_ sg13g2_and2_1
X_19772_ _12429_ VPWR VGND _12430_ sg13g2_buf_1
X_19773_ _08569_ _12430_ VPWR VGND _12431_ sg13g2_xnor2_1
X_19774_ _12399_ _12431_ VPWR VGND _12432_ sg13g2_nand2_1
X_19775_ _09106_ _12399_ _12432_ VPWR VGND _12433_ sg13g2_o21ai_1
X_19776_ \atbs_core_0.encoded_spike[12]\ _12394_ VPWR VGND _12434_ sg13g2_nand2_1
X_19777_ _12412_ _12433_ _12434_ VPWR VGND _00727_ sg13g2_o21ai_1
X_19778_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[13]\ VPWR VGND _12435_ sg13g2_buf_1
X_19779_ _12416_ _12420_ _12428_ VPWR VGND _12436_ sg13g2_nand3_1
X_19780_ _12436_ VPWR VGND _12437_ sg13g2_buf_1
X_19781_ _08854_ _12437_ VPWR VGND _12438_ sg13g2_nor2_1
X_19782_ _12435_ _12438_ VPWR VGND _12439_ sg13g2_xnor2_1
X_19783_ _09229_ _12424_ VPWR VGND _12440_ sg13g2_nor2_1
X_19784_ _12414_ _12439_ _12440_ VPWR VGND _12441_ sg13g2_a21oi_1
X_19785_ \atbs_core_0.encoded_spike[13]\ _12394_ VPWR VGND _12442_ sg13g2_nand2_1
X_19786_ _12412_ _12441_ _12442_ VPWR VGND _00728_ sg13g2_o21ai_1
X_19787_ _12435_ VPWR VGND _12443_ sg13g2_inv_1
X_19788_ _08569_ _12443_ _12430_ VPWR VGND _12444_ sg13g2_nand3_1
X_19789_ _09868_ _12444_ VPWR VGND _12445_ sg13g2_xnor2_1
X_19790_ _09720_ _12424_ VPWR VGND _12446_ sg13g2_nor2_1
X_19791_ _12414_ _12445_ _12446_ VPWR VGND _12447_ sg13g2_a21oi_1
X_19792_ \atbs_core_0.encoded_spike[14]\ _12394_ VPWR VGND _12448_ sg13g2_nand2_1
X_19793_ _12412_ _12447_ _12448_ VPWR VGND _00729_ sg13g2_o21ai_1
X_19794_ \atbs_core_0.adaptive_ctrl_0.curr_time_i[15]\ VPWR VGND _12449_ sg13g2_buf_1
X_19795_ _08943_ _08854_ _12435_ _12437_ VPWR VGND 
+ _12450_
+ sg13g2_nor4_1
X_19796_ _12449_ _12450_ VPWR VGND _12451_ sg13g2_xnor2_1
X_19797_ _08681_ _12424_ VPWR VGND _12452_ sg13g2_nor2_1
X_19798_ _12414_ _12451_ _12452_ VPWR VGND _12453_ sg13g2_a21oi_1
X_19799_ \atbs_core_0.encoded_spike[15]\ _12394_ VPWR VGND _12454_ sg13g2_nand2_1
X_19800_ _12412_ _12453_ _12454_ VPWR VGND _00730_ sg13g2_o21ai_1
X_19801_ _08684_ _08854_ _12435_ _12449_ VPWR VGND 
+ _12455_
+ sg13g2_nor4_1
X_19802_ _12430_ _12455_ VPWR VGND _12456_ sg13g2_nand2_1
X_19803_ _09035_ _12456_ VPWR VGND _12457_ sg13g2_xnor2_1
X_19804_ _08702_ _12424_ VPWR VGND _12458_ sg13g2_nor2_1
X_19805_ _12414_ _12457_ _12458_ VPWR VGND _12459_ sg13g2_a21oi_1
X_19806_ \atbs_core_0.encoded_spike[16]\ _12394_ VPWR VGND _12460_ sg13g2_nand2_1
X_19807_ _12412_ _12459_ _12460_ VPWR VGND _00731_ sg13g2_o21ai_1
X_19808_ _09035_ _12455_ VPWR VGND _12461_ sg13g2_and2_1
X_19809_ _12437_ _12461_ VPWR VGND _12462_ sg13g2_nor2b_1
X_19810_ _08709_ _12462_ VPWR VGND _12463_ sg13g2_xnor2_1
X_19811_ _08742_ _12424_ VPWR VGND _12464_ sg13g2_nor2_1
X_19812_ _12414_ _12463_ _12464_ VPWR VGND _12465_ sg13g2_a21oi_1
X_19813_ _12393_ VPWR VGND _12466_ sg13g2_buf_1
X_19814_ \atbs_core_0.encoded_spike[17]\ _12466_ VPWR VGND _12467_ sg13g2_nand2_1
X_19815_ _12412_ _12465_ _12467_ VPWR VGND _00732_ sg13g2_o21ai_1
X_19816_ _08762_ _12430_ _12461_ VPWR VGND _12468_ sg13g2_nand3_1
X_19817_ _07930_ _12414_ _12468_ VPWR VGND _12469_ sg13g2_nand3_1
X_19818_ \atbs_core_0.encoded_spike[18]\ _12466_ VPWR VGND _12470_ sg13g2_nand2_1
X_19819_ _12394_ _12469_ _12470_ VPWR VGND _00733_ sg13g2_o21ai_1
X_19820_ _08894_ _08892_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[1]\ sg13g2_xor2_1
X_19821_ _00023_ _12424_ VPWR VGND _12471_ sg13g2_nor2_1
X_19822_ _12414_ \atbs_core_0.time_measurement_0.n2218_o[1]\ _12471_ VPWR VGND _12472_ sg13g2_a21oi_1
X_19823_ \atbs_core_0.encoded_spike[1]\ _12466_ VPWR VGND _12473_ sg13g2_nand2_1
X_19824_ _12412_ _12472_ _12473_ VPWR VGND _00734_ sg13g2_o21ai_1
X_19825_ _08894_ _08892_ VPWR VGND _12474_ sg13g2_nor2_1
X_19826_ _08888_ _12474_ VPWR VGND _12475_ sg13g2_xnor2_1
X_19827_ _00024_ _12424_ VPWR VGND _12476_ sg13g2_nor2_1
X_19828_ _12414_ _12475_ _12476_ VPWR VGND _12477_ sg13g2_a21oi_1
X_19829_ \atbs_core_0.encoded_spike[2]\ _12466_ VPWR VGND _12478_ sg13g2_nand2_1
X_19830_ _12412_ _12477_ _12478_ VPWR VGND _00735_ sg13g2_o21ai_1
X_19831_ _08888_ _12417_ _08885_ VPWR VGND _12479_ sg13g2_o21ai_1
X_19832_ _12419_ _12479_ VPWR VGND _12480_ sg13g2_and2_1
X_19833_ _00025_ _12424_ VPWR VGND _12481_ sg13g2_nor2_1
X_19834_ _12414_ _12480_ _12481_ VPWR VGND _12482_ sg13g2_a21oi_1
X_19835_ \atbs_core_0.encoded_spike[3]\ _12466_ VPWR VGND _12483_ sg13g2_nand2_1
X_19836_ _12411_ _12482_ _12483_ VPWR VGND _00736_ sg13g2_o21ai_1
X_19837_ _08883_ _12401_ VPWR VGND _12484_ sg13g2_xnor2_1
X_19838_ _00026_ _12398_ VPWR VGND _12485_ sg13g2_nor2_1
X_19839_ _12399_ _12484_ _12485_ VPWR VGND _12486_ sg13g2_a21oi_1
X_19840_ \atbs_core_0.encoded_spike[4]\ _12466_ VPWR VGND _12487_ sg13g2_nand2_1
X_19841_ _12411_ _12486_ _12487_ VPWR VGND _00737_ sg13g2_o21ai_1
X_19842_ _08883_ _12419_ VPWR VGND _12488_ sg13g2_nor2_1
X_19843_ _08879_ _12488_ VPWR VGND _12489_ sg13g2_xnor2_1
X_19844_ _00027_ _12398_ VPWR VGND _12490_ sg13g2_nor2_1
X_19845_ _12399_ _12489_ _12490_ VPWR VGND _12491_ sg13g2_a21oi_1
X_19846_ \atbs_core_0.encoded_spike[5]\ _12466_ VPWR VGND _12492_ sg13g2_nand2_1
X_19847_ _12411_ _12491_ _12492_ VPWR VGND _00738_ sg13g2_o21ai_1
X_19848_ _08879_ _12402_ VPWR VGND _12493_ sg13g2_nor2_1
X_19849_ _08907_ _12493_ VPWR VGND _12494_ sg13g2_xnor2_1
X_19850_ _12399_ _12494_ VPWR VGND _12495_ sg13g2_nand2_1
X_19851_ _08475_ _12399_ _12495_ VPWR VGND _12496_ sg13g2_o21ai_1
X_19852_ \atbs_core_0.encoded_spike[6]\ _12466_ VPWR VGND _12497_ sg13g2_nand2_1
X_19853_ _12411_ _12496_ _12497_ VPWR VGND _00739_ sg13g2_o21ai_1
X_19854_ _12416_ _12420_ VPWR VGND _12498_ sg13g2_xnor2_1
X_19855_ _12424_ _12498_ VPWR VGND _12499_ sg13g2_nand2_1
X_19856_ _08534_ _12399_ _12499_ VPWR VGND _12500_ sg13g2_o21ai_1
X_19857_ \atbs_core_0.encoded_spike[7]\ _12466_ VPWR VGND _12501_ sg13g2_nand2_1
X_19858_ _12411_ _12500_ _12501_ VPWR VGND _00740_ sg13g2_o21ai_1
X_19859_ _10586_ _12403_ VPWR VGND _12502_ sg13g2_xnor2_1
X_19860_ _08549_ _12398_ VPWR VGND _12503_ sg13g2_nor2_1
X_19861_ _12399_ _12502_ _12503_ VPWR VGND _12504_ sg13g2_a21oi_1
X_19862_ \atbs_core_0.encoded_spike[8]\ _12466_ VPWR VGND _12505_ sg13g2_nand2_1
X_19863_ _12411_ _12504_ _12505_ VPWR VGND _00741_ sg13g2_o21ai_1
X_19864_ _10586_ _12421_ VPWR VGND _12506_ sg13g2_nor2_1
X_19865_ _12404_ _12506_ VPWR VGND _12507_ sg13g2_xnor2_1
X_19866_ _08577_ _12398_ VPWR VGND _12508_ sg13g2_nor2_1
X_19867_ _12399_ _12507_ _12508_ VPWR VGND _12509_ sg13g2_a21oi_1
X_19868_ \atbs_core_0.encoded_spike[9]\ _12393_ VPWR VGND _12510_ sg13g2_nand2_1
X_19869_ _12411_ _12509_ _12510_ VPWR VGND _00742_ sg13g2_o21ai_1
X_19870_ \atbs_core_0.spike_memory_0.n2439_q\ VPWR VGND _12511_ sg13g2_buf_1
X_19871_ _12511_ VPWR VGND _12512_ sg13g2_buf_1
X_19872_ _12512_ VPWR VGND _12513_ sg13g2_buf_1
X_19873_ _12513_ VPWR VGND _12514_ sg13g2_buf_1
X_19874_ \atbs_core_0.spike_memory_0.n2358_o[0]\ \atbs_core_0.spike_memory_0.a_data[0]\ _12514_ VPWR VGND _00743_ sg13g2_mux2_1
X_19875_ \atbs_core_0.spike_memory_0.n2410_o[12]\ \atbs_core_0.spike_memory_0.n2409_o[12]\ _12514_ VPWR VGND _00744_ sg13g2_mux2_1
X_19876_ \atbs_core_0.spike_memory_0.n2410_o[13]\ \atbs_core_0.spike_memory_0.n2409_o[13]\ _12514_ VPWR VGND _00745_ sg13g2_mux2_1
X_19877_ \atbs_core_0.spike_memory_0.n2410_o[14]\ \atbs_core_0.spike_memory_0.n2409_o[14]\ _12514_ VPWR VGND _00746_ sg13g2_mux2_1
X_19878_ \atbs_core_0.spike_memory_0.n2410_o[15]\ \atbs_core_0.spike_memory_0.n2409_o[15]\ _12514_ VPWR VGND _00747_ sg13g2_mux2_1
X_19879_ \atbs_core_0.spike_memory_0.n2410_o[16]\ \atbs_core_0.spike_memory_0.n2409_o[16]\ _12514_ VPWR VGND _00748_ sg13g2_mux2_1
X_19880_ _12513_ VPWR VGND _12515_ sg13g2_buf_1
X_19881_ \atbs_core_0.spike_memory_0.n2410_o[17]\ \atbs_core_0.spike_memory_0.n2409_o[17]\ _12515_ VPWR VGND _00749_ sg13g2_mux2_1
X_19882_ \atbs_core_0.spike_memory_0.n2410_o[18]\ \atbs_core_0.spike_memory_0.n2409_o[18]\ _12515_ VPWR VGND _00750_ sg13g2_mux2_1
X_19883_ \atbs_core_0.spike_memory_0.n2411_o[0]\ VPWR VGND _12516_ sg13g2_buf_1
X_19884_ _12516_ \atbs_core_0.spike_memory_0.n2410_o[0]\ _12515_ VPWR VGND _00751_ sg13g2_mux2_1
X_19885_ \atbs_core_0.spike_memory_0.n2411_o[1]\ VPWR VGND _12517_ sg13g2_buf_1
X_19886_ _12517_ \atbs_core_0.spike_memory_0.n2410_o[1]\ _12515_ VPWR VGND _00752_ sg13g2_mux2_1
X_19887_ \atbs_core_0.spike_memory_0.n2411_o[2]\ VPWR VGND _12518_ sg13g2_buf_1
X_19888_ _12518_ \atbs_core_0.spike_memory_0.n2410_o[2]\ _12515_ VPWR VGND _00753_ sg13g2_mux2_1
X_19889_ \atbs_core_0.spike_memory_0.n2363_o[5]\ VPWR VGND _12519_ sg13g2_buf_1
X_19890_ _12519_ \atbs_core_0.spike_memory_0.n2362_o[5]\ _12515_ VPWR VGND _00754_ sg13g2_mux2_1
X_19891_ \atbs_core_0.spike_memory_0.n2411_o[3]\ VPWR VGND _12520_ sg13g2_buf_1
X_19892_ _12520_ \atbs_core_0.spike_memory_0.n2410_o[3]\ _12515_ VPWR VGND _00755_ sg13g2_mux2_1
X_19893_ \atbs_core_0.spike_memory_0.n2411_o[4]\ VPWR VGND _12521_ sg13g2_buf_1
X_19894_ _12521_ \atbs_core_0.spike_memory_0.n2410_o[4]\ _12515_ VPWR VGND _00756_ sg13g2_mux2_1
X_19895_ \atbs_core_0.spike_memory_0.n2411_o[5]\ VPWR VGND _12522_ sg13g2_buf_1
X_19896_ _12522_ \atbs_core_0.spike_memory_0.n2410_o[5]\ _12515_ VPWR VGND _00757_ sg13g2_mux2_1
X_19897_ \atbs_core_0.spike_memory_0.n2411_o[6]\ VPWR VGND _12523_ sg13g2_buf_1
X_19898_ _12523_ \atbs_core_0.spike_memory_0.n2410_o[6]\ _12515_ VPWR VGND _00758_ sg13g2_mux2_1
X_19899_ \atbs_core_0.spike_memory_0.n2411_o[7]\ VPWR VGND _12524_ sg13g2_buf_1
X_19900_ _12512_ VPWR VGND _12525_ sg13g2_buf_1
X_19901_ _12525_ VPWR VGND _12526_ sg13g2_buf_1
X_19902_ _12524_ \atbs_core_0.spike_memory_0.n2410_o[7]\ _12526_ VPWR VGND _00759_ sg13g2_mux2_1
X_19903_ \atbs_core_0.spike_memory_0.n2411_o[8]\ VPWR VGND _12527_ sg13g2_buf_1
X_19904_ _12527_ \atbs_core_0.spike_memory_0.n2410_o[8]\ _12526_ VPWR VGND _00760_ sg13g2_mux2_1
X_19905_ \atbs_core_0.spike_memory_0.n2411_o[9]\ VPWR VGND _12528_ sg13g2_buf_1
X_19906_ _12528_ \atbs_core_0.spike_memory_0.n2410_o[9]\ _12526_ VPWR VGND _00761_ sg13g2_mux2_1
X_19907_ \atbs_core_0.spike_memory_0.n2411_o[10]\ VPWR VGND _12529_ sg13g2_buf_1
X_19908_ _12529_ \atbs_core_0.spike_memory_0.n2410_o[10]\ _12526_ VPWR VGND _00762_ sg13g2_mux2_1
X_19909_ \atbs_core_0.spike_memory_0.n2411_o[11]\ VPWR VGND _12530_ sg13g2_buf_1
X_19910_ _12530_ \atbs_core_0.spike_memory_0.n2410_o[11]\ _12526_ VPWR VGND _00763_ sg13g2_mux2_1
X_19911_ \atbs_core_0.spike_memory_0.n2411_o[12]\ VPWR VGND _12531_ sg13g2_buf_1
X_19912_ _12531_ \atbs_core_0.spike_memory_0.n2410_o[12]\ _12526_ VPWR VGND _00764_ sg13g2_mux2_1
X_19913_ \atbs_core_0.spike_memory_0.n2363_o[6]\ VPWR VGND _12532_ sg13g2_buf_1
X_19914_ _12532_ \atbs_core_0.spike_memory_0.n2362_o[6]\ _12526_ VPWR VGND _00765_ sg13g2_mux2_1
X_19915_ \atbs_core_0.spike_memory_0.n2411_o[13]\ VPWR VGND _12533_ sg13g2_buf_1
X_19916_ _12533_ \atbs_core_0.spike_memory_0.n2410_o[13]\ _12526_ VPWR VGND _00766_ sg13g2_mux2_1
X_19917_ \atbs_core_0.spike_memory_0.n2411_o[14]\ VPWR VGND _12534_ sg13g2_buf_1
X_19918_ _12534_ \atbs_core_0.spike_memory_0.n2410_o[14]\ _12526_ VPWR VGND _00767_ sg13g2_mux2_1
X_19919_ \atbs_core_0.spike_memory_0.n2411_o[15]\ VPWR VGND _12535_ sg13g2_buf_1
X_19920_ _12535_ \atbs_core_0.spike_memory_0.n2410_o[15]\ _12526_ VPWR VGND _00768_ sg13g2_mux2_1
X_19921_ \atbs_core_0.spike_memory_0.n2411_o[16]\ VPWR VGND _12536_ sg13g2_buf_1
X_19922_ _12525_ VPWR VGND _12537_ sg13g2_buf_1
X_19923_ _12536_ \atbs_core_0.spike_memory_0.n2410_o[16]\ _12537_ VPWR VGND _00769_ sg13g2_mux2_1
X_19924_ \atbs_core_0.spike_memory_0.n2411_o[17]\ VPWR VGND _12538_ sg13g2_buf_1
X_19925_ _12538_ \atbs_core_0.spike_memory_0.n2410_o[17]\ _12537_ VPWR VGND _00770_ sg13g2_mux2_1
X_19926_ \atbs_core_0.spike_memory_0.n2411_o[18]\ VPWR VGND _12539_ sg13g2_buf_1
X_19927_ _12539_ \atbs_core_0.spike_memory_0.n2410_o[18]\ _12537_ VPWR VGND _00771_ sg13g2_mux2_1
X_19928_ \atbs_core_0.spike_memory_0.n2412_o[0]\ VPWR VGND _12540_ sg13g2_buf_1
X_19929_ _12540_ _12516_ _12537_ VPWR VGND _00772_ sg13g2_mux2_1
X_19930_ \atbs_core_0.spike_memory_0.n2412_o[1]\ VPWR VGND _12541_ sg13g2_buf_1
X_19931_ _12541_ _12517_ _12537_ VPWR VGND _00773_ sg13g2_mux2_1
X_19932_ \atbs_core_0.spike_memory_0.n2412_o[2]\ VPWR VGND _12542_ sg13g2_buf_1
X_19933_ _12542_ _12518_ _12537_ VPWR VGND _00774_ sg13g2_mux2_1
X_19934_ \atbs_core_0.spike_memory_0.n2412_o[3]\ VPWR VGND _12543_ sg13g2_buf_1
X_19935_ _12543_ _12520_ _12537_ VPWR VGND _00775_ sg13g2_mux2_1
X_19936_ \atbs_core_0.spike_memory_0.n2363_o[7]\ VPWR VGND _12544_ sg13g2_buf_1
X_19937_ _12544_ \atbs_core_0.spike_memory_0.n2362_o[7]\ _12537_ VPWR VGND _00776_ sg13g2_mux2_1
X_19938_ \atbs_core_0.spike_memory_0.n2412_o[4]\ VPWR VGND _12545_ sg13g2_buf_1
X_19939_ _12545_ _12521_ _12537_ VPWR VGND _00777_ sg13g2_mux2_1
X_19940_ \atbs_core_0.spike_memory_0.n2412_o[5]\ VPWR VGND _12546_ sg13g2_buf_1
X_19941_ _12546_ _12522_ _12537_ VPWR VGND _00778_ sg13g2_mux2_1
X_19942_ \atbs_core_0.spike_memory_0.n2412_o[6]\ VPWR VGND _12547_ sg13g2_buf_1
X_19943_ _12525_ VPWR VGND _12548_ sg13g2_buf_1
X_19944_ _12547_ _12523_ _12548_ VPWR VGND _00779_ sg13g2_mux2_1
X_19945_ \atbs_core_0.spike_memory_0.n2412_o[7]\ VPWR VGND _12549_ sg13g2_buf_1
X_19946_ _12549_ _12524_ _12548_ VPWR VGND _00780_ sg13g2_mux2_1
X_19947_ \atbs_core_0.spike_memory_0.n2412_o[8]\ VPWR VGND _12550_ sg13g2_buf_1
X_19948_ _12550_ _12527_ _12548_ VPWR VGND _00781_ sg13g2_mux2_1
X_19949_ \atbs_core_0.spike_memory_0.n2412_o[9]\ VPWR VGND _12551_ sg13g2_buf_1
X_19950_ _12551_ _12528_ _12548_ VPWR VGND _00782_ sg13g2_mux2_1
X_19951_ \atbs_core_0.spike_memory_0.n2412_o[10]\ VPWR VGND _12552_ sg13g2_buf_1
X_19952_ _12552_ _12529_ _12548_ VPWR VGND _00783_ sg13g2_mux2_1
X_19953_ \atbs_core_0.spike_memory_0.n2412_o[11]\ VPWR VGND _12553_ sg13g2_buf_1
X_19954_ _12553_ _12530_ _12548_ VPWR VGND _00784_ sg13g2_mux2_1
X_19955_ \atbs_core_0.spike_memory_0.n2412_o[12]\ VPWR VGND _12554_ sg13g2_buf_1
X_19956_ _12554_ _12531_ _12548_ VPWR VGND _00785_ sg13g2_mux2_1
X_19957_ \atbs_core_0.spike_memory_0.n2412_o[13]\ VPWR VGND _12555_ sg13g2_buf_1
X_19958_ _12555_ _12533_ _12548_ VPWR VGND _00786_ sg13g2_mux2_1
X_19959_ \atbs_core_0.spike_memory_0.n2363_o[8]\ VPWR VGND _12556_ sg13g2_buf_1
X_19960_ _12556_ \atbs_core_0.spike_memory_0.n2362_o[8]\ _12548_ VPWR VGND _00787_ sg13g2_mux2_1
X_19961_ \atbs_core_0.spike_memory_0.n2412_o[14]\ VPWR VGND _12557_ sg13g2_buf_1
X_19962_ _12557_ _12534_ _12548_ VPWR VGND _00788_ sg13g2_mux2_1
X_19963_ \atbs_core_0.spike_memory_0.n2412_o[15]\ VPWR VGND _12558_ sg13g2_buf_1
X_19964_ _12525_ VPWR VGND _12559_ sg13g2_buf_1
X_19965_ _12558_ _12535_ _12559_ VPWR VGND _00789_ sg13g2_mux2_1
X_19966_ \atbs_core_0.spike_memory_0.n2412_o[16]\ VPWR VGND _12560_ sg13g2_buf_1
X_19967_ _12560_ _12536_ _12559_ VPWR VGND _00790_ sg13g2_mux2_1
X_19968_ \atbs_core_0.spike_memory_0.n2412_o[17]\ VPWR VGND _12561_ sg13g2_buf_1
X_19969_ _12561_ _12538_ _12559_ VPWR VGND _00791_ sg13g2_mux2_1
X_19970_ \atbs_core_0.spike_memory_0.n2412_o[18]\ VPWR VGND _12562_ sg13g2_buf_1
X_19971_ _12562_ _12539_ _12559_ VPWR VGND _00792_ sg13g2_mux2_1
X_19972_ \atbs_core_0.spike_memory_0.n2413_o[0]\ _12540_ _12559_ VPWR VGND _00793_ sg13g2_mux2_1
X_19973_ \atbs_core_0.spike_memory_0.n2413_o[1]\ _12541_ _12559_ VPWR VGND _00794_ sg13g2_mux2_1
X_19974_ \atbs_core_0.spike_memory_0.n2413_o[2]\ _12542_ _12559_ VPWR VGND _00795_ sg13g2_mux2_1
X_19975_ \atbs_core_0.spike_memory_0.n2413_o[3]\ _12543_ _12559_ VPWR VGND _00796_ sg13g2_mux2_1
X_19976_ \atbs_core_0.spike_memory_0.n2413_o[4]\ _12545_ _12559_ VPWR VGND _00797_ sg13g2_mux2_1
X_19977_ \atbs_core_0.spike_memory_0.n2363_o[9]\ VPWR VGND _12563_ sg13g2_buf_1
X_19978_ _12563_ \atbs_core_0.spike_memory_0.n2362_o[9]\ _12559_ VPWR VGND _00798_ sg13g2_mux2_1
X_19979_ _12525_ VPWR VGND _12564_ sg13g2_buf_1
X_19980_ \atbs_core_0.spike_memory_0.n2413_o[5]\ _12546_ _12564_ VPWR VGND _00799_ sg13g2_mux2_1
X_19981_ \atbs_core_0.spike_memory_0.n2413_o[6]\ _12547_ _12564_ VPWR VGND _00800_ sg13g2_mux2_1
X_19982_ \atbs_core_0.spike_memory_0.n2413_o[7]\ _12549_ _12564_ VPWR VGND _00801_ sg13g2_mux2_1
X_19983_ \atbs_core_0.spike_memory_0.n2413_o[8]\ _12550_ _12564_ VPWR VGND _00802_ sg13g2_mux2_1
X_19984_ \atbs_core_0.spike_memory_0.n2413_o[9]\ _12551_ _12564_ VPWR VGND _00803_ sg13g2_mux2_1
X_19985_ \atbs_core_0.spike_memory_0.n2413_o[10]\ _12552_ _12564_ VPWR VGND _00804_ sg13g2_mux2_1
X_19986_ \atbs_core_0.spike_memory_0.n2413_o[11]\ _12553_ _12564_ VPWR VGND _00805_ sg13g2_mux2_1
X_19987_ \atbs_core_0.spike_memory_0.n2413_o[12]\ _12554_ _12564_ VPWR VGND _00806_ sg13g2_mux2_1
X_19988_ \atbs_core_0.spike_memory_0.n2413_o[13]\ _12555_ _12564_ VPWR VGND _00807_ sg13g2_mux2_1
X_19989_ \atbs_core_0.spike_memory_0.n2413_o[14]\ _12557_ _12564_ VPWR VGND _00808_ sg13g2_mux2_1
X_19990_ \atbs_core_0.spike_memory_0.n2363_o[10]\ VPWR VGND _12565_ sg13g2_buf_1
X_19991_ _12525_ VPWR VGND _12566_ sg13g2_buf_1
X_19992_ _12565_ \atbs_core_0.spike_memory_0.n2362_o[10]\ _12566_ VPWR VGND _00809_ sg13g2_mux2_1
X_19993_ \atbs_core_0.spike_memory_0.n2413_o[15]\ _12558_ _12566_ VPWR VGND _00810_ sg13g2_mux2_1
X_19994_ \atbs_core_0.spike_memory_0.n2413_o[16]\ _12560_ _12566_ VPWR VGND _00811_ sg13g2_mux2_1
X_19995_ \atbs_core_0.spike_memory_0.n2413_o[17]\ _12561_ _12566_ VPWR VGND _00812_ sg13g2_mux2_1
X_19996_ \atbs_core_0.spike_memory_0.n2413_o[18]\ _12562_ _12566_ VPWR VGND _00813_ sg13g2_mux2_1
X_19997_ \atbs_core_0.spike_memory_0.n2414_o[0]\ \atbs_core_0.spike_memory_0.n2413_o[0]\ _12566_ VPWR VGND _00814_ sg13g2_mux2_1
X_19998_ \atbs_core_0.spike_memory_0.n2414_o[1]\ \atbs_core_0.spike_memory_0.n2413_o[1]\ _12566_ VPWR VGND _00815_ sg13g2_mux2_1
X_19999_ \atbs_core_0.spike_memory_0.n2414_o[2]\ \atbs_core_0.spike_memory_0.n2413_o[2]\ _12566_ VPWR VGND _00816_ sg13g2_mux2_1
X_20000_ \atbs_core_0.spike_memory_0.n2414_o[3]\ \atbs_core_0.spike_memory_0.n2413_o[3]\ _12566_ VPWR VGND _00817_ sg13g2_mux2_1
X_20001_ \atbs_core_0.spike_memory_0.n2414_o[4]\ \atbs_core_0.spike_memory_0.n2413_o[4]\ _12566_ VPWR VGND _00818_ sg13g2_mux2_1
X_20002_ _12525_ VPWR VGND _12567_ sg13g2_buf_1
X_20003_ \atbs_core_0.spike_memory_0.n2414_o[5]\ \atbs_core_0.spike_memory_0.n2413_o[5]\ _12567_ VPWR VGND _00819_ sg13g2_mux2_1
X_20004_ \atbs_core_0.spike_memory_0.n2363_o[11]\ VPWR VGND _12568_ sg13g2_buf_1
X_20005_ _12568_ \atbs_core_0.spike_memory_0.n2362_o[11]\ _12567_ VPWR VGND _00820_ sg13g2_mux2_1
X_20006_ \atbs_core_0.spike_memory_0.n2414_o[6]\ \atbs_core_0.spike_memory_0.n2413_o[6]\ _12567_ VPWR VGND _00821_ sg13g2_mux2_1
X_20007_ \atbs_core_0.spike_memory_0.n2414_o[7]\ \atbs_core_0.spike_memory_0.n2413_o[7]\ _12567_ VPWR VGND _00822_ sg13g2_mux2_1
X_20008_ \atbs_core_0.spike_memory_0.n2414_o[8]\ \atbs_core_0.spike_memory_0.n2413_o[8]\ _12567_ VPWR VGND _00823_ sg13g2_mux2_1
X_20009_ \atbs_core_0.spike_memory_0.n2414_o[9]\ \atbs_core_0.spike_memory_0.n2413_o[9]\ _12567_ VPWR VGND _00824_ sg13g2_mux2_1
X_20010_ \atbs_core_0.spike_memory_0.n2414_o[10]\ \atbs_core_0.spike_memory_0.n2413_o[10]\ _12567_ VPWR VGND _00825_ sg13g2_mux2_1
X_20011_ \atbs_core_0.spike_memory_0.n2414_o[11]\ \atbs_core_0.spike_memory_0.n2413_o[11]\ _12567_ VPWR VGND _00826_ sg13g2_mux2_1
X_20012_ \atbs_core_0.spike_memory_0.n2414_o[12]\ \atbs_core_0.spike_memory_0.n2413_o[12]\ _12567_ VPWR VGND _00827_ sg13g2_mux2_1
X_20013_ \atbs_core_0.spike_memory_0.n2414_o[13]\ \atbs_core_0.spike_memory_0.n2413_o[13]\ _12567_ VPWR VGND _00828_ sg13g2_mux2_1
X_20014_ _12512_ VPWR VGND _12569_ sg13g2_buf_1
X_20015_ _12569_ VPWR VGND _12570_ sg13g2_buf_1
X_20016_ \atbs_core_0.spike_memory_0.n2414_o[14]\ \atbs_core_0.spike_memory_0.n2413_o[14]\ _12570_ VPWR VGND _00829_ sg13g2_mux2_1
X_20017_ \atbs_core_0.spike_memory_0.n2414_o[15]\ \atbs_core_0.spike_memory_0.n2413_o[15]\ _12570_ VPWR VGND _00830_ sg13g2_mux2_1
X_20018_ \atbs_core_0.spike_memory_0.n2363_o[12]\ VPWR VGND _12571_ sg13g2_buf_1
X_20019_ _12571_ \atbs_core_0.spike_memory_0.n2362_o[12]\ _12570_ VPWR VGND _00831_ sg13g2_mux2_1
X_20020_ \atbs_core_0.spike_memory_0.n2414_o[16]\ \atbs_core_0.spike_memory_0.n2413_o[16]\ _12570_ VPWR VGND _00832_ sg13g2_mux2_1
X_20021_ \atbs_core_0.spike_memory_0.n2414_o[17]\ \atbs_core_0.spike_memory_0.n2413_o[17]\ _12570_ VPWR VGND _00833_ sg13g2_mux2_1
X_20022_ \atbs_core_0.spike_memory_0.n2414_o[18]\ \atbs_core_0.spike_memory_0.n2413_o[18]\ _12570_ VPWR VGND _00834_ sg13g2_mux2_1
X_20023_ \atbs_core_0.spike_memory_0.n2415_o[0]\ VPWR VGND _12572_ sg13g2_buf_1
X_20024_ _12572_ \atbs_core_0.spike_memory_0.n2414_o[0]\ _12570_ VPWR VGND _00835_ sg13g2_mux2_1
X_20025_ \atbs_core_0.spike_memory_0.n2415_o[1]\ VPWR VGND _12573_ sg13g2_buf_1
X_20026_ _12573_ \atbs_core_0.spike_memory_0.n2414_o[1]\ _12570_ VPWR VGND _00836_ sg13g2_mux2_1
X_20027_ \atbs_core_0.spike_memory_0.n2415_o[2]\ VPWR VGND _12574_ sg13g2_buf_1
X_20028_ _12574_ \atbs_core_0.spike_memory_0.n2414_o[2]\ _12570_ VPWR VGND _00837_ sg13g2_mux2_1
X_20029_ \atbs_core_0.spike_memory_0.n2415_o[3]\ VPWR VGND _12575_ sg13g2_buf_1
X_20030_ _12575_ \atbs_core_0.spike_memory_0.n2414_o[3]\ _12570_ VPWR VGND _00838_ sg13g2_mux2_1
X_20031_ \atbs_core_0.spike_memory_0.n2415_o[4]\ VPWR VGND _12576_ sg13g2_buf_1
X_20032_ _12569_ VPWR VGND _12577_ sg13g2_buf_1
X_20033_ _12576_ \atbs_core_0.spike_memory_0.n2414_o[4]\ _12577_ VPWR VGND _00839_ sg13g2_mux2_1
X_20034_ \atbs_core_0.spike_memory_0.n2415_o[5]\ VPWR VGND _12578_ sg13g2_buf_1
X_20035_ _12578_ \atbs_core_0.spike_memory_0.n2414_o[5]\ _12577_ VPWR VGND _00840_ sg13g2_mux2_1
X_20036_ \atbs_core_0.spike_memory_0.n2415_o[6]\ VPWR VGND _12579_ sg13g2_buf_1
X_20037_ _12579_ \atbs_core_0.spike_memory_0.n2414_o[6]\ _12577_ VPWR VGND _00841_ sg13g2_mux2_1
X_20038_ \atbs_core_0.spike_memory_0.n2363_o[13]\ VPWR VGND _12580_ sg13g2_buf_1
X_20039_ _12580_ \atbs_core_0.spike_memory_0.n2362_o[13]\ _12577_ VPWR VGND _00842_ sg13g2_mux2_1
X_20040_ \atbs_core_0.spike_memory_0.n2415_o[7]\ VPWR VGND _12581_ sg13g2_buf_1
X_20041_ _12581_ \atbs_core_0.spike_memory_0.n2414_o[7]\ _12577_ VPWR VGND _00843_ sg13g2_mux2_1
X_20042_ \atbs_core_0.spike_memory_0.n2415_o[8]\ VPWR VGND _12582_ sg13g2_buf_1
X_20043_ _12582_ \atbs_core_0.spike_memory_0.n2414_o[8]\ _12577_ VPWR VGND _00844_ sg13g2_mux2_1
X_20044_ \atbs_core_0.spike_memory_0.n2415_o[9]\ VPWR VGND _12583_ sg13g2_buf_1
X_20045_ _12583_ \atbs_core_0.spike_memory_0.n2414_o[9]\ _12577_ VPWR VGND _00845_ sg13g2_mux2_1
X_20046_ \atbs_core_0.spike_memory_0.n2415_o[10]\ VPWR VGND _12584_ sg13g2_buf_1
X_20047_ _12584_ \atbs_core_0.spike_memory_0.n2414_o[10]\ _12577_ VPWR VGND _00846_ sg13g2_mux2_1
X_20048_ \atbs_core_0.spike_memory_0.n2415_o[11]\ VPWR VGND _12585_ sg13g2_buf_1
X_20049_ _12585_ \atbs_core_0.spike_memory_0.n2414_o[11]\ _12577_ VPWR VGND _00847_ sg13g2_mux2_1
X_20050_ \atbs_core_0.spike_memory_0.n2415_o[12]\ VPWR VGND _12586_ sg13g2_buf_1
X_20051_ _12586_ \atbs_core_0.spike_memory_0.n2414_o[12]\ _12577_ VPWR VGND _00848_ sg13g2_mux2_1
X_20052_ \atbs_core_0.spike_memory_0.n2415_o[13]\ VPWR VGND _12587_ sg13g2_buf_1
X_20053_ _12569_ VPWR VGND _12588_ sg13g2_buf_1
X_20054_ _12587_ \atbs_core_0.spike_memory_0.n2414_o[13]\ _12588_ VPWR VGND _00849_ sg13g2_mux2_1
X_20055_ \atbs_core_0.spike_memory_0.n2415_o[14]\ VPWR VGND _12589_ sg13g2_buf_1
X_20056_ _12589_ \atbs_core_0.spike_memory_0.n2414_o[14]\ _12588_ VPWR VGND _00850_ sg13g2_mux2_1
X_20057_ \atbs_core_0.spike_memory_0.n2415_o[15]\ VPWR VGND _12590_ sg13g2_buf_1
X_20058_ _12590_ \atbs_core_0.spike_memory_0.n2414_o[15]\ _12588_ VPWR VGND _00851_ sg13g2_mux2_1
X_20059_ \atbs_core_0.spike_memory_0.n2415_o[16]\ VPWR VGND _12591_ sg13g2_buf_1
X_20060_ _12591_ \atbs_core_0.spike_memory_0.n2414_o[16]\ _12588_ VPWR VGND _00852_ sg13g2_mux2_1
X_20061_ \atbs_core_0.spike_memory_0.n2363_o[14]\ VPWR VGND _12592_ sg13g2_buf_1
X_20062_ _12592_ \atbs_core_0.spike_memory_0.n2362_o[14]\ _12588_ VPWR VGND _00853_ sg13g2_mux2_1
X_20063_ \atbs_core_0.spike_memory_0.n2358_o[10]\ \atbs_core_0.spike_memory_0.a_data[10]\ _12588_ VPWR VGND _00854_ sg13g2_mux2_1
X_20064_ \atbs_core_0.spike_memory_0.n2415_o[17]\ VPWR VGND _12593_ sg13g2_buf_1
X_20065_ _12593_ \atbs_core_0.spike_memory_0.n2414_o[17]\ _12588_ VPWR VGND _00855_ sg13g2_mux2_1
X_20066_ \atbs_core_0.spike_memory_0.n2415_o[18]\ VPWR VGND _12594_ sg13g2_buf_1
X_20067_ _12594_ \atbs_core_0.spike_memory_0.n2414_o[18]\ _12588_ VPWR VGND _00856_ sg13g2_mux2_1
X_20068_ \atbs_core_0.spike_memory_0.n2416_o[0]\ VPWR VGND _12595_ sg13g2_buf_1
X_20069_ _12595_ _12572_ _12588_ VPWR VGND _00857_ sg13g2_mux2_1
X_20070_ \atbs_core_0.spike_memory_0.n2416_o[1]\ VPWR VGND _12596_ sg13g2_buf_1
X_20071_ _12596_ _12573_ _12588_ VPWR VGND _00858_ sg13g2_mux2_1
X_20072_ \atbs_core_0.spike_memory_0.n2416_o[2]\ VPWR VGND _12597_ sg13g2_buf_1
X_20073_ _12569_ VPWR VGND _12598_ sg13g2_buf_1
X_20074_ _12597_ _12574_ _12598_ VPWR VGND _00859_ sg13g2_mux2_1
X_20075_ \atbs_core_0.spike_memory_0.n2416_o[3]\ VPWR VGND _12599_ sg13g2_buf_1
X_20076_ _12599_ _12575_ _12598_ VPWR VGND _00860_ sg13g2_mux2_1
X_20077_ \atbs_core_0.spike_memory_0.n2416_o[4]\ VPWR VGND _12600_ sg13g2_buf_1
X_20078_ _12600_ _12576_ _12598_ VPWR VGND _00861_ sg13g2_mux2_1
X_20079_ \atbs_core_0.spike_memory_0.n2416_o[5]\ VPWR VGND _12601_ sg13g2_buf_1
X_20080_ _12601_ _12578_ _12598_ VPWR VGND _00862_ sg13g2_mux2_1
X_20081_ \atbs_core_0.spike_memory_0.n2416_o[6]\ VPWR VGND _12602_ sg13g2_buf_1
X_20082_ _12602_ _12579_ _12598_ VPWR VGND _00863_ sg13g2_mux2_1
X_20083_ \atbs_core_0.spike_memory_0.n2416_o[7]\ VPWR VGND _12603_ sg13g2_buf_1
X_20084_ _12603_ _12581_ _12598_ VPWR VGND _00864_ sg13g2_mux2_1
X_20085_ \atbs_core_0.spike_memory_0.n2363_o[15]\ VPWR VGND _12604_ sg13g2_buf_1
X_20086_ _12604_ \atbs_core_0.spike_memory_0.n2362_o[15]\ _12598_ VPWR VGND _00865_ sg13g2_mux2_1
X_20087_ \atbs_core_0.spike_memory_0.n2416_o[8]\ VPWR VGND _12605_ sg13g2_buf_1
X_20088_ _12605_ _12582_ _12598_ VPWR VGND _00866_ sg13g2_mux2_1
X_20089_ \atbs_core_0.spike_memory_0.n2416_o[9]\ VPWR VGND _12606_ sg13g2_buf_1
X_20090_ _12606_ _12583_ _12598_ VPWR VGND _00867_ sg13g2_mux2_1
X_20091_ \atbs_core_0.spike_memory_0.n2416_o[10]\ VPWR VGND _12607_ sg13g2_buf_1
X_20092_ _12607_ _12584_ _12598_ VPWR VGND _00868_ sg13g2_mux2_1
X_20093_ \atbs_core_0.spike_memory_0.n2416_o[11]\ VPWR VGND _12608_ sg13g2_buf_1
X_20094_ _12569_ VPWR VGND _12609_ sg13g2_buf_1
X_20095_ _12608_ _12585_ _12609_ VPWR VGND _00869_ sg13g2_mux2_1
X_20096_ \atbs_core_0.spike_memory_0.n2416_o[12]\ VPWR VGND _12610_ sg13g2_buf_1
X_20097_ _12610_ _12586_ _12609_ VPWR VGND _00870_ sg13g2_mux2_1
X_20098_ \atbs_core_0.spike_memory_0.n2416_o[13]\ VPWR VGND _12611_ sg13g2_buf_1
X_20099_ _12611_ _12587_ _12609_ VPWR VGND _00871_ sg13g2_mux2_1
X_20100_ \atbs_core_0.spike_memory_0.n2416_o[14]\ VPWR VGND _12612_ sg13g2_buf_1
X_20101_ _12612_ _12589_ _12609_ VPWR VGND _00872_ sg13g2_mux2_1
X_20102_ \atbs_core_0.spike_memory_0.n2416_o[15]\ VPWR VGND _12613_ sg13g2_buf_1
X_20103_ _12613_ _12590_ _12609_ VPWR VGND _00873_ sg13g2_mux2_1
X_20104_ \atbs_core_0.spike_memory_0.n2416_o[16]\ VPWR VGND _12614_ sg13g2_buf_1
X_20105_ _12614_ _12591_ _12609_ VPWR VGND _00874_ sg13g2_mux2_1
X_20106_ \atbs_core_0.spike_memory_0.n2416_o[17]\ VPWR VGND _12615_ sg13g2_buf_1
X_20107_ _12615_ _12593_ _12609_ VPWR VGND _00875_ sg13g2_mux2_1
X_20108_ \atbs_core_0.spike_memory_0.n2363_o[16]\ VPWR VGND _12616_ sg13g2_buf_1
X_20109_ _12616_ \atbs_core_0.spike_memory_0.n2362_o[16]\ _12609_ VPWR VGND _00876_ sg13g2_mux2_1
X_20110_ \atbs_core_0.spike_memory_0.n2416_o[18]\ VPWR VGND _12617_ sg13g2_buf_1
X_20111_ _12617_ _12594_ _12609_ VPWR VGND _00877_ sg13g2_mux2_1
X_20112_ \atbs_core_0.spike_memory_0.n2417_o[0]\ _12595_ _12609_ VPWR VGND _00878_ sg13g2_mux2_1
X_20113_ _12569_ VPWR VGND _12618_ sg13g2_buf_1
X_20114_ \atbs_core_0.spike_memory_0.n2417_o[1]\ _12596_ _12618_ VPWR VGND _00879_ sg13g2_mux2_1
X_20115_ \atbs_core_0.spike_memory_0.n2417_o[2]\ _12597_ _12618_ VPWR VGND _00880_ sg13g2_mux2_1
X_20116_ \atbs_core_0.spike_memory_0.n2417_o[3]\ _12599_ _12618_ VPWR VGND _00881_ sg13g2_mux2_1
X_20117_ \atbs_core_0.spike_memory_0.n2417_o[4]\ _12600_ _12618_ VPWR VGND _00882_ sg13g2_mux2_1
X_20118_ \atbs_core_0.spike_memory_0.n2417_o[5]\ _12601_ _12618_ VPWR VGND _00883_ sg13g2_mux2_1
X_20119_ \atbs_core_0.spike_memory_0.n2417_o[6]\ _12602_ _12618_ VPWR VGND _00884_ sg13g2_mux2_1
X_20120_ \atbs_core_0.spike_memory_0.n2417_o[7]\ _12603_ _12618_ VPWR VGND _00885_ sg13g2_mux2_1
X_20121_ \atbs_core_0.spike_memory_0.n2417_o[8]\ _12605_ _12618_ VPWR VGND _00886_ sg13g2_mux2_1
X_20122_ \atbs_core_0.spike_memory_0.n2363_o[17]\ VPWR VGND _12619_ sg13g2_buf_1
X_20123_ _12619_ \atbs_core_0.spike_memory_0.n2362_o[17]\ _12618_ VPWR VGND _00887_ sg13g2_mux2_1
X_20124_ \atbs_core_0.spike_memory_0.n2417_o[9]\ _12606_ _12618_ VPWR VGND _00888_ sg13g2_mux2_1
X_20125_ _12569_ VPWR VGND _12620_ sg13g2_buf_1
X_20126_ \atbs_core_0.spike_memory_0.n2417_o[10]\ _12607_ _12620_ VPWR VGND _00889_ sg13g2_mux2_1
X_20127_ \atbs_core_0.spike_memory_0.n2417_o[11]\ _12608_ _12620_ VPWR VGND _00890_ sg13g2_mux2_1
X_20128_ \atbs_core_0.spike_memory_0.n2417_o[12]\ _12610_ _12620_ VPWR VGND _00891_ sg13g2_mux2_1
X_20129_ \atbs_core_0.spike_memory_0.n2417_o[13]\ _12611_ _12620_ VPWR VGND _00892_ sg13g2_mux2_1
X_20130_ \atbs_core_0.spike_memory_0.n2417_o[14]\ _12612_ _12620_ VPWR VGND _00893_ sg13g2_mux2_1
X_20131_ \atbs_core_0.spike_memory_0.n2417_o[15]\ _12613_ _12620_ VPWR VGND _00894_ sg13g2_mux2_1
X_20132_ \atbs_core_0.spike_memory_0.n2417_o[16]\ _12614_ _12620_ VPWR VGND _00895_ sg13g2_mux2_1
X_20133_ \atbs_core_0.spike_memory_0.n2417_o[17]\ _12615_ _12620_ VPWR VGND _00896_ sg13g2_mux2_1
X_20134_ \atbs_core_0.spike_memory_0.n2417_o[18]\ _12617_ _12620_ VPWR VGND _00897_ sg13g2_mux2_1
X_20135_ \atbs_core_0.spike_memory_0.n2363_o[18]\ VPWR VGND _12621_ sg13g2_buf_1
X_20136_ _12621_ \atbs_core_0.spike_memory_0.n2362_o[18]\ _12620_ VPWR VGND _00898_ sg13g2_mux2_1
X_20137_ _12512_ VPWR VGND _12622_ sg13g2_buf_1
X_20138_ _12622_ VPWR VGND _12623_ sg13g2_buf_1
X_20139_ \atbs_core_0.spike_memory_0.n2418_o[0]\ \atbs_core_0.spike_memory_0.n2417_o[0]\ _12623_ VPWR VGND _00899_ sg13g2_mux2_1
X_20140_ \atbs_core_0.spike_memory_0.n2418_o[1]\ \atbs_core_0.spike_memory_0.n2417_o[1]\ _12623_ VPWR VGND _00900_ sg13g2_mux2_1
X_20141_ \atbs_core_0.spike_memory_0.n2418_o[2]\ \atbs_core_0.spike_memory_0.n2417_o[2]\ _12623_ VPWR VGND _00901_ sg13g2_mux2_1
X_20142_ \atbs_core_0.spike_memory_0.n2418_o[3]\ \atbs_core_0.spike_memory_0.n2417_o[3]\ _12623_ VPWR VGND _00902_ sg13g2_mux2_1
X_20143_ \atbs_core_0.spike_memory_0.n2418_o[4]\ \atbs_core_0.spike_memory_0.n2417_o[4]\ _12623_ VPWR VGND _00903_ sg13g2_mux2_1
X_20144_ \atbs_core_0.spike_memory_0.n2418_o[5]\ \atbs_core_0.spike_memory_0.n2417_o[5]\ _12623_ VPWR VGND _00904_ sg13g2_mux2_1
X_20145_ \atbs_core_0.spike_memory_0.n2418_o[6]\ \atbs_core_0.spike_memory_0.n2417_o[6]\ _12623_ VPWR VGND _00905_ sg13g2_mux2_1
X_20146_ \atbs_core_0.spike_memory_0.n2418_o[7]\ \atbs_core_0.spike_memory_0.n2417_o[7]\ _12623_ VPWR VGND _00906_ sg13g2_mux2_1
X_20147_ \atbs_core_0.spike_memory_0.n2418_o[8]\ \atbs_core_0.spike_memory_0.n2417_o[8]\ _12623_ VPWR VGND _00907_ sg13g2_mux2_1
X_20148_ \atbs_core_0.spike_memory_0.n2418_o[9]\ \atbs_core_0.spike_memory_0.n2417_o[9]\ _12623_ VPWR VGND _00908_ sg13g2_mux2_1
X_20149_ \atbs_core_0.spike_memory_0.n2364_o[0]\ VPWR VGND _12624_ sg13g2_buf_1
X_20150_ \atbs_core_0.spike_memory_0.n2363_o[0]\ VPWR VGND _12625_ sg13g2_buf_1
X_20151_ _12622_ VPWR VGND _12626_ sg13g2_buf_1
X_20152_ _12624_ _12625_ _12626_ VPWR VGND _00909_ sg13g2_mux2_1
X_20153_ \atbs_core_0.spike_memory_0.n2418_o[10]\ \atbs_core_0.spike_memory_0.n2417_o[10]\ _12626_ VPWR VGND _00910_ sg13g2_mux2_1
X_20154_ \atbs_core_0.spike_memory_0.n2418_o[11]\ \atbs_core_0.spike_memory_0.n2417_o[11]\ _12626_ VPWR VGND _00911_ sg13g2_mux2_1
X_20155_ \atbs_core_0.spike_memory_0.n2418_o[12]\ \atbs_core_0.spike_memory_0.n2417_o[12]\ _12626_ VPWR VGND _00912_ sg13g2_mux2_1
X_20156_ \atbs_core_0.spike_memory_0.n2418_o[13]\ \atbs_core_0.spike_memory_0.n2417_o[13]\ _12626_ VPWR VGND _00913_ sg13g2_mux2_1
X_20157_ \atbs_core_0.spike_memory_0.n2418_o[14]\ \atbs_core_0.spike_memory_0.n2417_o[14]\ _12626_ VPWR VGND _00914_ sg13g2_mux2_1
X_20158_ \atbs_core_0.spike_memory_0.n2418_o[15]\ \atbs_core_0.spike_memory_0.n2417_o[15]\ _12626_ VPWR VGND _00915_ sg13g2_mux2_1
X_20159_ \atbs_core_0.spike_memory_0.n2418_o[16]\ \atbs_core_0.spike_memory_0.n2417_o[16]\ _12626_ VPWR VGND _00916_ sg13g2_mux2_1
X_20160_ \atbs_core_0.spike_memory_0.n2418_o[17]\ \atbs_core_0.spike_memory_0.n2417_o[17]\ _12626_ VPWR VGND _00917_ sg13g2_mux2_1
X_20161_ \atbs_core_0.spike_memory_0.n2418_o[18]\ \atbs_core_0.spike_memory_0.n2417_o[18]\ _12626_ VPWR VGND _00918_ sg13g2_mux2_1
X_20162_ \atbs_core_0.spike_memory_0.n2419_o[0]\ VPWR VGND _12627_ sg13g2_buf_1
X_20163_ _12622_ VPWR VGND _12628_ sg13g2_buf_1
X_20164_ _12627_ \atbs_core_0.spike_memory_0.n2418_o[0]\ _12628_ VPWR VGND _00919_ sg13g2_mux2_1
X_20165_ \atbs_core_0.spike_memory_0.n2364_o[1]\ VPWR VGND _12629_ sg13g2_buf_1
X_20166_ \atbs_core_0.spike_memory_0.n2363_o[1]\ VPWR VGND _12630_ sg13g2_buf_1
X_20167_ _12629_ _12630_ _12628_ VPWR VGND _00920_ sg13g2_mux2_1
X_20168_ \atbs_core_0.spike_memory_0.n2419_o[1]\ VPWR VGND _12631_ sg13g2_buf_1
X_20169_ _12631_ \atbs_core_0.spike_memory_0.n2418_o[1]\ _12628_ VPWR VGND _00921_ sg13g2_mux2_1
X_20170_ \atbs_core_0.spike_memory_0.n2419_o[2]\ VPWR VGND _12632_ sg13g2_buf_1
X_20171_ _12632_ \atbs_core_0.spike_memory_0.n2418_o[2]\ _12628_ VPWR VGND _00922_ sg13g2_mux2_1
X_20172_ \atbs_core_0.spike_memory_0.n2419_o[3]\ VPWR VGND _12633_ sg13g2_buf_1
X_20173_ _12633_ \atbs_core_0.spike_memory_0.n2418_o[3]\ _12628_ VPWR VGND _00923_ sg13g2_mux2_1
X_20174_ \atbs_core_0.spike_memory_0.n2419_o[4]\ VPWR VGND _12634_ sg13g2_buf_1
X_20175_ _12634_ \atbs_core_0.spike_memory_0.n2418_o[4]\ _12628_ VPWR VGND _00924_ sg13g2_mux2_1
X_20176_ \atbs_core_0.spike_memory_0.n2419_o[5]\ VPWR VGND _12635_ sg13g2_buf_1
X_20177_ _12635_ \atbs_core_0.spike_memory_0.n2418_o[5]\ _12628_ VPWR VGND _00925_ sg13g2_mux2_1
X_20178_ \atbs_core_0.spike_memory_0.n2419_o[6]\ VPWR VGND _12636_ sg13g2_buf_1
X_20179_ _12636_ \atbs_core_0.spike_memory_0.n2418_o[6]\ _12628_ VPWR VGND _00926_ sg13g2_mux2_1
X_20180_ \atbs_core_0.spike_memory_0.n2419_o[7]\ VPWR VGND _12637_ sg13g2_buf_1
X_20181_ _12637_ \atbs_core_0.spike_memory_0.n2418_o[7]\ _12628_ VPWR VGND _00927_ sg13g2_mux2_1
X_20182_ \atbs_core_0.spike_memory_0.n2419_o[8]\ VPWR VGND _12638_ sg13g2_buf_1
X_20183_ _12638_ \atbs_core_0.spike_memory_0.n2418_o[8]\ _12628_ VPWR VGND _00928_ sg13g2_mux2_1
X_20184_ \atbs_core_0.spike_memory_0.n2419_o[9]\ VPWR VGND _12639_ sg13g2_buf_1
X_20185_ _12622_ VPWR VGND _12640_ sg13g2_buf_1
X_20186_ _12639_ \atbs_core_0.spike_memory_0.n2418_o[9]\ _12640_ VPWR VGND _00929_ sg13g2_mux2_1
X_20187_ \atbs_core_0.spike_memory_0.n2419_o[10]\ VPWR VGND _12641_ sg13g2_buf_1
X_20188_ _12641_ \atbs_core_0.spike_memory_0.n2418_o[10]\ _12640_ VPWR VGND _00930_ sg13g2_mux2_1
X_20189_ \atbs_core_0.spike_memory_0.n2364_o[2]\ VPWR VGND _12642_ sg13g2_buf_1
X_20190_ \atbs_core_0.spike_memory_0.n2363_o[2]\ VPWR VGND _12643_ sg13g2_buf_1
X_20191_ _12642_ _12643_ _12640_ VPWR VGND _00931_ sg13g2_mux2_1
X_20192_ \atbs_core_0.spike_memory_0.n2419_o[11]\ VPWR VGND _12644_ sg13g2_buf_1
X_20193_ _12644_ \atbs_core_0.spike_memory_0.n2418_o[11]\ _12640_ VPWR VGND _00932_ sg13g2_mux2_1
X_20194_ \atbs_core_0.spike_memory_0.n2419_o[12]\ VPWR VGND _12645_ sg13g2_buf_1
X_20195_ _12645_ \atbs_core_0.spike_memory_0.n2418_o[12]\ _12640_ VPWR VGND _00933_ sg13g2_mux2_1
X_20196_ \atbs_core_0.spike_memory_0.n2419_o[13]\ VPWR VGND _12646_ sg13g2_buf_1
X_20197_ _12646_ \atbs_core_0.spike_memory_0.n2418_o[13]\ _12640_ VPWR VGND _00934_ sg13g2_mux2_1
X_20198_ \atbs_core_0.spike_memory_0.n2419_o[14]\ VPWR VGND _12647_ sg13g2_buf_1
X_20199_ _12647_ \atbs_core_0.spike_memory_0.n2418_o[14]\ _12640_ VPWR VGND _00935_ sg13g2_mux2_1
X_20200_ \atbs_core_0.spike_memory_0.n2419_o[15]\ VPWR VGND _12648_ sg13g2_buf_1
X_20201_ _12648_ \atbs_core_0.spike_memory_0.n2418_o[15]\ _12640_ VPWR VGND _00936_ sg13g2_mux2_1
X_20202_ \atbs_core_0.spike_memory_0.n2419_o[16]\ VPWR VGND _12649_ sg13g2_buf_1
X_20203_ _12649_ \atbs_core_0.spike_memory_0.n2418_o[16]\ _12640_ VPWR VGND _00937_ sg13g2_mux2_1
X_20204_ \atbs_core_0.spike_memory_0.n2419_o[17]\ VPWR VGND _12650_ sg13g2_buf_1
X_20205_ _12650_ \atbs_core_0.spike_memory_0.n2418_o[17]\ _12640_ VPWR VGND _00938_ sg13g2_mux2_1
X_20206_ \atbs_core_0.spike_memory_0.n2419_o[18]\ VPWR VGND _12651_ sg13g2_buf_1
X_20207_ _12622_ VPWR VGND _12652_ sg13g2_buf_1
X_20208_ _12651_ \atbs_core_0.spike_memory_0.n2418_o[18]\ _12652_ VPWR VGND _00939_ sg13g2_mux2_1
X_20209_ \atbs_core_0.spike_memory_0.n2420_o[0]\ VPWR VGND _12653_ sg13g2_buf_1
X_20210_ _12653_ _12627_ _12652_ VPWR VGND _00940_ sg13g2_mux2_1
X_20211_ \atbs_core_0.spike_memory_0.n2420_o[1]\ VPWR VGND _12654_ sg13g2_buf_1
X_20212_ _12654_ _12631_ _12652_ VPWR VGND _00941_ sg13g2_mux2_1
X_20213_ \atbs_core_0.spike_memory_0.n2364_o[3]\ VPWR VGND _12655_ sg13g2_buf_1
X_20214_ \atbs_core_0.spike_memory_0.n2363_o[3]\ VPWR VGND _12656_ sg13g2_buf_1
X_20215_ _12655_ _12656_ _12652_ VPWR VGND _00942_ sg13g2_mux2_1
X_20216_ \atbs_core_0.spike_memory_0.n2420_o[2]\ VPWR VGND _12657_ sg13g2_buf_1
X_20217_ _12657_ _12632_ _12652_ VPWR VGND _00943_ sg13g2_mux2_1
X_20218_ \atbs_core_0.spike_memory_0.n2420_o[3]\ VPWR VGND _12658_ sg13g2_buf_1
X_20219_ _12658_ _12633_ _12652_ VPWR VGND _00944_ sg13g2_mux2_1
X_20220_ \atbs_core_0.spike_memory_0.n2420_o[4]\ VPWR VGND _12659_ sg13g2_buf_1
X_20221_ _12659_ _12634_ _12652_ VPWR VGND _00945_ sg13g2_mux2_1
X_20222_ \atbs_core_0.spike_memory_0.n2420_o[5]\ VPWR VGND _12660_ sg13g2_buf_1
X_20223_ _12660_ _12635_ _12652_ VPWR VGND _00946_ sg13g2_mux2_1
X_20224_ \atbs_core_0.spike_memory_0.n2420_o[6]\ VPWR VGND _12661_ sg13g2_buf_1
X_20225_ _12661_ _12636_ _12652_ VPWR VGND _00947_ sg13g2_mux2_1
X_20226_ \atbs_core_0.spike_memory_0.n2420_o[7]\ VPWR VGND _12662_ sg13g2_buf_1
X_20227_ _12662_ _12637_ _12652_ VPWR VGND _00948_ sg13g2_mux2_1
X_20228_ \atbs_core_0.spike_memory_0.n2420_o[8]\ VPWR VGND _12663_ sg13g2_buf_1
X_20229_ _12622_ VPWR VGND _12664_ sg13g2_buf_1
X_20230_ _12663_ _12638_ _12664_ VPWR VGND _00949_ sg13g2_mux2_1
X_20231_ \atbs_core_0.spike_memory_0.n2420_o[9]\ VPWR VGND _12665_ sg13g2_buf_1
X_20232_ _12665_ _12639_ _12664_ VPWR VGND _00950_ sg13g2_mux2_1
X_20233_ \atbs_core_0.spike_memory_0.n2420_o[10]\ VPWR VGND _12666_ sg13g2_buf_1
X_20234_ _12666_ _12641_ _12664_ VPWR VGND _00951_ sg13g2_mux2_1
X_20235_ \atbs_core_0.spike_memory_0.n2420_o[11]\ VPWR VGND _12667_ sg13g2_buf_1
X_20236_ _12667_ _12644_ _12664_ VPWR VGND _00952_ sg13g2_mux2_1
X_20237_ \atbs_core_0.spike_memory_0.n2364_o[4]\ VPWR VGND _12668_ sg13g2_buf_1
X_20238_ \atbs_core_0.spike_memory_0.n2363_o[4]\ VPWR VGND _12669_ sg13g2_buf_1
X_20239_ _12668_ _12669_ _12664_ VPWR VGND _00953_ sg13g2_mux2_1
X_20240_ \atbs_core_0.spike_memory_0.n2420_o[12]\ VPWR VGND _12670_ sg13g2_buf_1
X_20241_ _12670_ _12645_ _12664_ VPWR VGND _00954_ sg13g2_mux2_1
X_20242_ \atbs_core_0.spike_memory_0.n2420_o[13]\ VPWR VGND _12671_ sg13g2_buf_1
X_20243_ _12671_ _12646_ _12664_ VPWR VGND _00955_ sg13g2_mux2_1
X_20244_ \atbs_core_0.spike_memory_0.n2420_o[14]\ VPWR VGND _12672_ sg13g2_buf_1
X_20245_ _12672_ _12647_ _12664_ VPWR VGND _00956_ sg13g2_mux2_1
X_20246_ \atbs_core_0.spike_memory_0.n2420_o[15]\ VPWR VGND _12673_ sg13g2_buf_1
X_20247_ _12673_ _12648_ _12664_ VPWR VGND _00957_ sg13g2_mux2_1
X_20248_ \atbs_core_0.spike_memory_0.n2420_o[16]\ VPWR VGND _12674_ sg13g2_buf_1
X_20249_ _12674_ _12649_ _12664_ VPWR VGND _00958_ sg13g2_mux2_1
X_20250_ \atbs_core_0.spike_memory_0.n2420_o[17]\ VPWR VGND _12675_ sg13g2_buf_1
X_20251_ _12622_ VPWR VGND _12676_ sg13g2_buf_1
X_20252_ _12675_ _12650_ _12676_ VPWR VGND _00959_ sg13g2_mux2_1
X_20253_ \atbs_core_0.spike_memory_0.n2420_o[18]\ VPWR VGND _12677_ sg13g2_buf_1
X_20254_ _12677_ _12651_ _12676_ VPWR VGND _00960_ sg13g2_mux2_1
X_20255_ \atbs_core_0.spike_memory_0.n2436_q[1197]\ _12653_ _12676_ VPWR VGND _00961_ sg13g2_mux2_1
X_20256_ \atbs_core_0.spike_memory_0.n2436_q[1198]\ _12654_ _12676_ VPWR VGND _00962_ sg13g2_mux2_1
X_20257_ \atbs_core_0.spike_memory_0.n2436_q[1199]\ _12657_ _12676_ VPWR VGND _00963_ sg13g2_mux2_1
X_20258_ \atbs_core_0.spike_memory_0.n2364_o[5]\ VPWR VGND _12678_ sg13g2_buf_1
X_20259_ _12678_ _12519_ _12676_ VPWR VGND _00964_ sg13g2_mux2_1
X_20260_ \atbs_core_0.spike_memory_0.n2358_o[11]\ \atbs_core_0.spike_memory_0.a_data[11]\ _12676_ VPWR VGND _00965_ sg13g2_mux2_1
X_20261_ \atbs_core_0.spike_memory_0.n2436_q[1200]\ _12658_ _12676_ VPWR VGND _00966_ sg13g2_mux2_1
X_20262_ \atbs_core_0.spike_memory_0.n2436_q[1201]\ _12659_ _12676_ VPWR VGND _00967_ sg13g2_mux2_1
X_20263_ \atbs_core_0.spike_memory_0.n2436_q[1202]\ _12660_ _12676_ VPWR VGND _00968_ sg13g2_mux2_1
X_20264_ _12512_ VPWR VGND _12679_ sg13g2_buf_1
X_20265_ _12679_ VPWR VGND _12680_ sg13g2_buf_1
X_20266_ \atbs_core_0.spike_memory_0.n2436_q[1203]\ _12661_ _12680_ VPWR VGND _00969_ sg13g2_mux2_1
X_20267_ \atbs_core_0.spike_memory_0.n2436_q[1204]\ _12662_ _12680_ VPWR VGND _00970_ sg13g2_mux2_1
X_20268_ \atbs_core_0.spike_memory_0.n2436_q[1205]\ _12663_ _12680_ VPWR VGND _00971_ sg13g2_mux2_1
X_20269_ \atbs_core_0.spike_memory_0.n2436_q[1206]\ _12665_ _12680_ VPWR VGND _00972_ sg13g2_mux2_1
X_20270_ \atbs_core_0.spike_memory_0.n2436_q[1207]\ _12666_ _12680_ VPWR VGND _00973_ sg13g2_mux2_1
X_20271_ \atbs_core_0.spike_memory_0.n2436_q[1208]\ _12667_ _12680_ VPWR VGND _00974_ sg13g2_mux2_1
X_20272_ \atbs_core_0.spike_memory_0.n2436_q[1209]\ _12670_ _12680_ VPWR VGND _00975_ sg13g2_mux2_1
X_20273_ \atbs_core_0.spike_memory_0.n2364_o[6]\ VPWR VGND _12681_ sg13g2_buf_1
X_20274_ _12681_ _12532_ _12680_ VPWR VGND _00976_ sg13g2_mux2_1
X_20275_ \atbs_core_0.spike_memory_0.n2436_q[1210]\ _12671_ _12680_ VPWR VGND _00977_ sg13g2_mux2_1
X_20276_ \atbs_core_0.spike_memory_0.n2436_q[1211]\ _12672_ _12680_ VPWR VGND _00978_ sg13g2_mux2_1
X_20277_ _12679_ VPWR VGND _12682_ sg13g2_buf_1
X_20278_ \atbs_core_0.spike_memory_0.n2436_q[1212]\ _12673_ _12682_ VPWR VGND _00979_ sg13g2_mux2_1
X_20279_ \atbs_core_0.spike_memory_0.n2436_q[1213]\ _12674_ _12682_ VPWR VGND _00980_ sg13g2_mux2_1
X_20280_ \atbs_core_0.spike_memory_0.n2436_q[1214]\ _12675_ _12682_ VPWR VGND _00981_ sg13g2_mux2_1
X_20281_ \atbs_core_0.spike_memory_0.n2436_q[1215]\ _12677_ _12682_ VPWR VGND _00982_ sg13g2_mux2_1
X_20282_ \atbs_core_0.spike_memory_0.n2364_o[7]\ VPWR VGND _02007_ sg13g2_buf_1
X_20283_ _02007_ _12544_ _12682_ VPWR VGND _00983_ sg13g2_mux2_1
X_20284_ \atbs_core_0.spike_memory_0.n2364_o[8]\ VPWR VGND _02008_ sg13g2_buf_1
X_20285_ _02008_ _12556_ _12682_ VPWR VGND _00984_ sg13g2_mux2_1
X_20286_ \atbs_core_0.spike_memory_0.n2364_o[9]\ VPWR VGND _02009_ sg13g2_buf_1
X_20287_ _02009_ _12563_ _12682_ VPWR VGND _00985_ sg13g2_mux2_1
X_20288_ \atbs_core_0.spike_memory_0.n2364_o[10]\ VPWR VGND _02010_ sg13g2_buf_1
X_20289_ _02010_ _12565_ _12682_ VPWR VGND _00986_ sg13g2_mux2_1
X_20290_ \atbs_core_0.spike_memory_0.n2364_o[11]\ VPWR VGND _02011_ sg13g2_buf_1
X_20291_ _02011_ _12568_ _12682_ VPWR VGND _00987_ sg13g2_mux2_1
X_20292_ \atbs_core_0.spike_memory_0.n2364_o[12]\ VPWR VGND _02012_ sg13g2_buf_1
X_20293_ _02012_ _12571_ _12682_ VPWR VGND _00988_ sg13g2_mux2_1
X_20294_ \atbs_core_0.spike_memory_0.n2364_o[13]\ VPWR VGND _02013_ sg13g2_buf_1
X_20295_ _12679_ VPWR VGND _02014_ sg13g2_buf_1
X_20296_ _02013_ _12580_ _02014_ VPWR VGND _00989_ sg13g2_mux2_1
X_20297_ \atbs_core_0.spike_memory_0.n2364_o[14]\ VPWR VGND _02015_ sg13g2_buf_1
X_20298_ _02015_ _12592_ _02014_ VPWR VGND _00990_ sg13g2_mux2_1
X_20299_ \atbs_core_0.spike_memory_0.n2364_o[15]\ VPWR VGND _02016_ sg13g2_buf_1
X_20300_ _02016_ _12604_ _02014_ VPWR VGND _00991_ sg13g2_mux2_1
X_20301_ \atbs_core_0.spike_memory_0.n2358_o[12]\ \atbs_core_0.spike_memory_0.a_data[12]\ _02014_ VPWR VGND _00992_ sg13g2_mux2_1
X_20302_ \atbs_core_0.spike_memory_0.n2364_o[16]\ VPWR VGND _02017_ sg13g2_buf_1
X_20303_ _02017_ _12616_ _02014_ VPWR VGND _00993_ sg13g2_mux2_1
X_20304_ \atbs_core_0.spike_memory_0.n2364_o[17]\ VPWR VGND _02018_ sg13g2_buf_1
X_20305_ _02018_ _12619_ _02014_ VPWR VGND _00994_ sg13g2_mux2_1
X_20306_ \atbs_core_0.spike_memory_0.n2364_o[18]\ VPWR VGND _02019_ sg13g2_buf_1
X_20307_ _02019_ _12621_ _02014_ VPWR VGND _00995_ sg13g2_mux2_1
X_20308_ \atbs_core_0.spike_memory_0.n2365_o[0]\ _12624_ _02014_ VPWR VGND _00996_ sg13g2_mux2_1
X_20309_ \atbs_core_0.spike_memory_0.n2365_o[1]\ _12629_ _02014_ VPWR VGND _00997_ sg13g2_mux2_1
X_20310_ \atbs_core_0.spike_memory_0.n2365_o[2]\ _12642_ _02014_ VPWR VGND _00998_ sg13g2_mux2_1
X_20311_ _12679_ VPWR VGND _02020_ sg13g2_buf_1
X_20312_ \atbs_core_0.spike_memory_0.n2365_o[3]\ _12655_ _02020_ VPWR VGND _00999_ sg13g2_mux2_1
X_20313_ \atbs_core_0.spike_memory_0.n2365_o[4]\ _12668_ _02020_ VPWR VGND _01000_ sg13g2_mux2_1
X_20314_ \atbs_core_0.spike_memory_0.n2365_o[5]\ _12678_ _02020_ VPWR VGND _01001_ sg13g2_mux2_1
X_20315_ \atbs_core_0.spike_memory_0.n2365_o[6]\ _12681_ _02020_ VPWR VGND _01002_ sg13g2_mux2_1
X_20316_ \atbs_core_0.spike_memory_0.n2358_o[13]\ \atbs_core_0.spike_memory_0.a_data[13]\ _02020_ VPWR VGND _01003_ sg13g2_mux2_1
X_20317_ \atbs_core_0.spike_memory_0.n2365_o[7]\ _02007_ _02020_ VPWR VGND _01004_ sg13g2_mux2_1
X_20318_ \atbs_core_0.spike_memory_0.n2365_o[8]\ _02008_ _02020_ VPWR VGND _01005_ sg13g2_mux2_1
X_20319_ \atbs_core_0.spike_memory_0.n2365_o[9]\ _02009_ _02020_ VPWR VGND _01006_ sg13g2_mux2_1
X_20320_ \atbs_core_0.spike_memory_0.n2365_o[10]\ _02010_ _02020_ VPWR VGND _01007_ sg13g2_mux2_1
X_20321_ \atbs_core_0.spike_memory_0.n2365_o[11]\ _02011_ _02020_ VPWR VGND _01008_ sg13g2_mux2_1
X_20322_ _12679_ VPWR VGND _02021_ sg13g2_buf_1
X_20323_ \atbs_core_0.spike_memory_0.n2365_o[12]\ _02012_ _02021_ VPWR VGND _01009_ sg13g2_mux2_1
X_20324_ \atbs_core_0.spike_memory_0.n2365_o[13]\ _02013_ _02021_ VPWR VGND _01010_ sg13g2_mux2_1
X_20325_ \atbs_core_0.spike_memory_0.n2365_o[14]\ _02015_ _02021_ VPWR VGND _01011_ sg13g2_mux2_1
X_20326_ \atbs_core_0.spike_memory_0.n2365_o[15]\ _02016_ _02021_ VPWR VGND _01012_ sg13g2_mux2_1
X_20327_ \atbs_core_0.spike_memory_0.n2365_o[16]\ _02017_ _02021_ VPWR VGND _01013_ sg13g2_mux2_1
X_20328_ \atbs_core_0.spike_memory_0.n2358_o[14]\ \atbs_core_0.spike_memory_0.a_data[14]\ _02021_ VPWR VGND _01014_ sg13g2_mux2_1
X_20329_ \atbs_core_0.spike_memory_0.n2365_o[17]\ _02018_ _02021_ VPWR VGND _01015_ sg13g2_mux2_1
X_20330_ \atbs_core_0.spike_memory_0.n2365_o[18]\ _02019_ _02021_ VPWR VGND _01016_ sg13g2_mux2_1
X_20331_ \atbs_core_0.spike_memory_0.n2366_o[0]\ \atbs_core_0.spike_memory_0.n2365_o[0]\ _02021_ VPWR VGND _01017_ sg13g2_mux2_1
X_20332_ \atbs_core_0.spike_memory_0.n2366_o[1]\ \atbs_core_0.spike_memory_0.n2365_o[1]\ _02021_ VPWR VGND _01018_ sg13g2_mux2_1
X_20333_ _12679_ VPWR VGND _02022_ sg13g2_buf_1
X_20334_ \atbs_core_0.spike_memory_0.n2366_o[2]\ \atbs_core_0.spike_memory_0.n2365_o[2]\ _02022_ VPWR VGND _01019_ sg13g2_mux2_1
X_20335_ \atbs_core_0.spike_memory_0.n2366_o[3]\ \atbs_core_0.spike_memory_0.n2365_o[3]\ _02022_ VPWR VGND _01020_ sg13g2_mux2_1
X_20336_ \atbs_core_0.spike_memory_0.n2366_o[4]\ \atbs_core_0.spike_memory_0.n2365_o[4]\ _02022_ VPWR VGND _01021_ sg13g2_mux2_1
X_20337_ \atbs_core_0.spike_memory_0.n2366_o[5]\ \atbs_core_0.spike_memory_0.n2365_o[5]\ _02022_ VPWR VGND _01022_ sg13g2_mux2_1
X_20338_ \atbs_core_0.spike_memory_0.n2366_o[6]\ \atbs_core_0.spike_memory_0.n2365_o[6]\ _02022_ VPWR VGND _01023_ sg13g2_mux2_1
X_20339_ \atbs_core_0.spike_memory_0.n2366_o[7]\ \atbs_core_0.spike_memory_0.n2365_o[7]\ _02022_ VPWR VGND _01024_ sg13g2_mux2_1
X_20340_ \atbs_core_0.spike_memory_0.n2358_o[15]\ \atbs_core_0.spike_memory_0.a_data[15]\ _02022_ VPWR VGND _01025_ sg13g2_mux2_1
X_20341_ \atbs_core_0.spike_memory_0.n2366_o[8]\ \atbs_core_0.spike_memory_0.n2365_o[8]\ _02022_ VPWR VGND _01026_ sg13g2_mux2_1
X_20342_ \atbs_core_0.spike_memory_0.n2366_o[9]\ \atbs_core_0.spike_memory_0.n2365_o[9]\ _02022_ VPWR VGND _01027_ sg13g2_mux2_1
X_20343_ \atbs_core_0.spike_memory_0.n2366_o[10]\ \atbs_core_0.spike_memory_0.n2365_o[10]\ _02022_ VPWR VGND _01028_ sg13g2_mux2_1
X_20344_ _12679_ VPWR VGND _02023_ sg13g2_buf_1
X_20345_ \atbs_core_0.spike_memory_0.n2366_o[11]\ \atbs_core_0.spike_memory_0.n2365_o[11]\ _02023_ VPWR VGND _01029_ sg13g2_mux2_1
X_20346_ \atbs_core_0.spike_memory_0.n2366_o[12]\ \atbs_core_0.spike_memory_0.n2365_o[12]\ _02023_ VPWR VGND _01030_ sg13g2_mux2_1
X_20347_ \atbs_core_0.spike_memory_0.n2366_o[13]\ \atbs_core_0.spike_memory_0.n2365_o[13]\ _02023_ VPWR VGND _01031_ sg13g2_mux2_1
X_20348_ \atbs_core_0.spike_memory_0.n2366_o[14]\ \atbs_core_0.spike_memory_0.n2365_o[14]\ _02023_ VPWR VGND _01032_ sg13g2_mux2_1
X_20349_ \atbs_core_0.spike_memory_0.n2366_o[15]\ \atbs_core_0.spike_memory_0.n2365_o[15]\ _02023_ VPWR VGND _01033_ sg13g2_mux2_1
X_20350_ \atbs_core_0.spike_memory_0.n2366_o[16]\ \atbs_core_0.spike_memory_0.n2365_o[16]\ _02023_ VPWR VGND _01034_ sg13g2_mux2_1
X_20351_ \atbs_core_0.spike_memory_0.n2366_o[17]\ \atbs_core_0.spike_memory_0.n2365_o[17]\ _02023_ VPWR VGND _01035_ sg13g2_mux2_1
X_20352_ \atbs_core_0.spike_memory_0.n2358_o[16]\ \atbs_core_0.spike_memory_0.a_data[16]\ _02023_ VPWR VGND _01036_ sg13g2_mux2_1
X_20353_ \atbs_core_0.spike_memory_0.n2366_o[18]\ \atbs_core_0.spike_memory_0.n2365_o[18]\ _02023_ VPWR VGND _01037_ sg13g2_mux2_1
X_20354_ \atbs_core_0.spike_memory_0.n2367_o[0]\ VPWR VGND _02024_ sg13g2_buf_1
X_20355_ _02024_ \atbs_core_0.spike_memory_0.n2366_o[0]\ _02023_ VPWR VGND _01038_ sg13g2_mux2_1
X_20356_ \atbs_core_0.spike_memory_0.n2367_o[1]\ VPWR VGND _02025_ sg13g2_buf_1
X_20357_ _12512_ VPWR VGND _02026_ sg13g2_buf_1
X_20358_ _02026_ VPWR VGND _02027_ sg13g2_buf_1
X_20359_ _02025_ \atbs_core_0.spike_memory_0.n2366_o[1]\ _02027_ VPWR VGND _01039_ sg13g2_mux2_1
X_20360_ \atbs_core_0.spike_memory_0.n2367_o[2]\ VPWR VGND _02028_ sg13g2_buf_1
X_20361_ _02028_ \atbs_core_0.spike_memory_0.n2366_o[2]\ _02027_ VPWR VGND _01040_ sg13g2_mux2_1
X_20362_ \atbs_core_0.spike_memory_0.n2367_o[3]\ VPWR VGND _02029_ sg13g2_buf_1
X_20363_ _02029_ \atbs_core_0.spike_memory_0.n2366_o[3]\ _02027_ VPWR VGND _01041_ sg13g2_mux2_1
X_20364_ \atbs_core_0.spike_memory_0.n2367_o[4]\ VPWR VGND _02030_ sg13g2_buf_1
X_20365_ _02030_ \atbs_core_0.spike_memory_0.n2366_o[4]\ _02027_ VPWR VGND _01042_ sg13g2_mux2_1
X_20366_ \atbs_core_0.spike_memory_0.n2367_o[5]\ VPWR VGND _02031_ sg13g2_buf_1
X_20367_ _02031_ \atbs_core_0.spike_memory_0.n2366_o[5]\ _02027_ VPWR VGND _01043_ sg13g2_mux2_1
X_20368_ \atbs_core_0.spike_memory_0.n2367_o[6]\ VPWR VGND _02032_ sg13g2_buf_1
X_20369_ _02032_ \atbs_core_0.spike_memory_0.n2366_o[6]\ _02027_ VPWR VGND _01044_ sg13g2_mux2_1
X_20370_ \atbs_core_0.spike_memory_0.n2367_o[7]\ VPWR VGND _02033_ sg13g2_buf_1
X_20371_ _02033_ \atbs_core_0.spike_memory_0.n2366_o[7]\ _02027_ VPWR VGND _01045_ sg13g2_mux2_1
X_20372_ \atbs_core_0.spike_memory_0.n2367_o[8]\ VPWR VGND _02034_ sg13g2_buf_1
X_20373_ _02034_ \atbs_core_0.spike_memory_0.n2366_o[8]\ _02027_ VPWR VGND _01046_ sg13g2_mux2_1
X_20374_ \atbs_core_0.spike_memory_0.n2358_o[17]\ \atbs_core_0.spike_memory_0.a_data[17]\ _02027_ VPWR VGND _01047_ sg13g2_mux2_1
X_20375_ \atbs_core_0.spike_memory_0.n2367_o[9]\ VPWR VGND _02035_ sg13g2_buf_1
X_20376_ _02035_ \atbs_core_0.spike_memory_0.n2366_o[9]\ _02027_ VPWR VGND _01048_ sg13g2_mux2_1
X_20377_ \atbs_core_0.spike_memory_0.n2367_o[10]\ VPWR VGND _02036_ sg13g2_buf_1
X_20378_ _02026_ VPWR VGND _02037_ sg13g2_buf_1
X_20379_ _02036_ \atbs_core_0.spike_memory_0.n2366_o[10]\ _02037_ VPWR VGND _01049_ sg13g2_mux2_1
X_20380_ \atbs_core_0.spike_memory_0.n2367_o[11]\ VPWR VGND _02038_ sg13g2_buf_1
X_20381_ _02038_ \atbs_core_0.spike_memory_0.n2366_o[11]\ _02037_ VPWR VGND _01050_ sg13g2_mux2_1
X_20382_ \atbs_core_0.spike_memory_0.n2367_o[12]\ VPWR VGND _02039_ sg13g2_buf_1
X_20383_ _02039_ \atbs_core_0.spike_memory_0.n2366_o[12]\ _02037_ VPWR VGND _01051_ sg13g2_mux2_1
X_20384_ \atbs_core_0.spike_memory_0.n2367_o[13]\ VPWR VGND _02040_ sg13g2_buf_1
X_20385_ _02040_ \atbs_core_0.spike_memory_0.n2366_o[13]\ _02037_ VPWR VGND _01052_ sg13g2_mux2_1
X_20386_ \atbs_core_0.spike_memory_0.n2367_o[14]\ VPWR VGND _02041_ sg13g2_buf_1
X_20387_ _02041_ \atbs_core_0.spike_memory_0.n2366_o[14]\ _02037_ VPWR VGND _01053_ sg13g2_mux2_1
X_20388_ \atbs_core_0.spike_memory_0.n2367_o[15]\ VPWR VGND _02042_ sg13g2_buf_1
X_20389_ _02042_ \atbs_core_0.spike_memory_0.n2366_o[15]\ _02037_ VPWR VGND _01054_ sg13g2_mux2_1
X_20390_ \atbs_core_0.spike_memory_0.n2367_o[16]\ VPWR VGND _02043_ sg13g2_buf_1
X_20391_ _02043_ \atbs_core_0.spike_memory_0.n2366_o[16]\ _02037_ VPWR VGND _01055_ sg13g2_mux2_1
X_20392_ \atbs_core_0.spike_memory_0.n2367_o[17]\ VPWR VGND _02044_ sg13g2_buf_1
X_20393_ _02044_ \atbs_core_0.spike_memory_0.n2366_o[17]\ _02037_ VPWR VGND _01056_ sg13g2_mux2_1
X_20394_ \atbs_core_0.spike_memory_0.n2367_o[18]\ VPWR VGND _02045_ sg13g2_buf_1
X_20395_ _02045_ \atbs_core_0.spike_memory_0.n2366_o[18]\ _02037_ VPWR VGND _01057_ sg13g2_mux2_1
X_20396_ \atbs_core_0.spike_memory_0.n2358_o[18]\ \atbs_core_0.spike_memory_0.a_data[18]\ _02037_ VPWR VGND _01058_ sg13g2_mux2_1
X_20397_ \atbs_core_0.spike_memory_0.n2368_o[0]\ VPWR VGND _02046_ sg13g2_buf_1
X_20398_ _02026_ VPWR VGND _02047_ sg13g2_buf_1
X_20399_ _02046_ _02024_ _02047_ VPWR VGND _01059_ sg13g2_mux2_1
X_20400_ \atbs_core_0.spike_memory_0.n2368_o[1]\ VPWR VGND _02048_ sg13g2_buf_1
X_20401_ _02048_ _02025_ _02047_ VPWR VGND _01060_ sg13g2_mux2_1
X_20402_ \atbs_core_0.spike_memory_0.n2368_o[2]\ VPWR VGND _02049_ sg13g2_buf_1
X_20403_ _02049_ _02028_ _02047_ VPWR VGND _01061_ sg13g2_mux2_1
X_20404_ \atbs_core_0.spike_memory_0.n2368_o[3]\ VPWR VGND _02050_ sg13g2_buf_1
X_20405_ _02050_ _02029_ _02047_ VPWR VGND _01062_ sg13g2_mux2_1
X_20406_ \atbs_core_0.spike_memory_0.n2368_o[4]\ VPWR VGND _02051_ sg13g2_buf_1
X_20407_ _02051_ _02030_ _02047_ VPWR VGND _01063_ sg13g2_mux2_1
X_20408_ \atbs_core_0.spike_memory_0.n2368_o[5]\ VPWR VGND _02052_ sg13g2_buf_1
X_20409_ _02052_ _02031_ _02047_ VPWR VGND _01064_ sg13g2_mux2_1
X_20410_ \atbs_core_0.spike_memory_0.n2368_o[6]\ VPWR VGND _02053_ sg13g2_buf_1
X_20411_ _02053_ _02032_ _02047_ VPWR VGND _01065_ sg13g2_mux2_1
X_20412_ \atbs_core_0.spike_memory_0.n2368_o[7]\ VPWR VGND _02054_ sg13g2_buf_1
X_20413_ _02054_ _02033_ _02047_ VPWR VGND _01066_ sg13g2_mux2_1
X_20414_ \atbs_core_0.spike_memory_0.n2368_o[8]\ VPWR VGND _02055_ sg13g2_buf_1
X_20415_ _02055_ _02034_ _02047_ VPWR VGND _01067_ sg13g2_mux2_1
X_20416_ \atbs_core_0.spike_memory_0.n2368_o[9]\ VPWR VGND _02056_ sg13g2_buf_1
X_20417_ _02056_ _02035_ _02047_ VPWR VGND _01068_ sg13g2_mux2_1
X_20418_ \atbs_core_0.spike_memory_0.n2359_o[0]\ VPWR VGND _02057_ sg13g2_buf_1
X_20419_ _02026_ VPWR VGND _02058_ sg13g2_buf_1
X_20420_ _02057_ \atbs_core_0.spike_memory_0.n2358_o[0]\ _02058_ VPWR VGND _01069_ sg13g2_mux2_1
X_20421_ \atbs_core_0.spike_memory_0.n2358_o[1]\ \atbs_core_0.spike_memory_0.a_data[1]\ _02058_ VPWR VGND _01070_ sg13g2_mux2_1
X_20422_ \atbs_core_0.spike_memory_0.n2368_o[10]\ VPWR VGND _02059_ sg13g2_buf_1
X_20423_ _02059_ _02036_ _02058_ VPWR VGND _01071_ sg13g2_mux2_1
X_20424_ \atbs_core_0.spike_memory_0.n2368_o[11]\ VPWR VGND _02060_ sg13g2_buf_1
X_20425_ _02060_ _02038_ _02058_ VPWR VGND _01072_ sg13g2_mux2_1
X_20426_ \atbs_core_0.spike_memory_0.n2368_o[12]\ VPWR VGND _02061_ sg13g2_buf_1
X_20427_ _02061_ _02039_ _02058_ VPWR VGND _01073_ sg13g2_mux2_1
X_20428_ \atbs_core_0.spike_memory_0.n2368_o[13]\ VPWR VGND _02062_ sg13g2_buf_1
X_20429_ _02062_ _02040_ _02058_ VPWR VGND _01074_ sg13g2_mux2_1
X_20430_ \atbs_core_0.spike_memory_0.n2368_o[14]\ VPWR VGND _02063_ sg13g2_buf_1
X_20431_ _02063_ _02041_ _02058_ VPWR VGND _01075_ sg13g2_mux2_1
X_20432_ \atbs_core_0.spike_memory_0.n2368_o[15]\ VPWR VGND _02064_ sg13g2_buf_1
X_20433_ _02064_ _02042_ _02058_ VPWR VGND _01076_ sg13g2_mux2_1
X_20434_ \atbs_core_0.spike_memory_0.n2368_o[16]\ VPWR VGND _02065_ sg13g2_buf_1
X_20435_ _02065_ _02043_ _02058_ VPWR VGND _01077_ sg13g2_mux2_1
X_20436_ \atbs_core_0.spike_memory_0.n2368_o[17]\ VPWR VGND _02066_ sg13g2_buf_1
X_20437_ _02066_ _02044_ _02058_ VPWR VGND _01078_ sg13g2_mux2_1
X_20438_ \atbs_core_0.spike_memory_0.n2368_o[18]\ VPWR VGND _02067_ sg13g2_buf_1
X_20439_ _02026_ VPWR VGND _02068_ sg13g2_buf_1
X_20440_ _02067_ _02045_ _02068_ VPWR VGND _01079_ sg13g2_mux2_1
X_20441_ \atbs_core_0.spike_memory_0.n2369_o[0]\ _02046_ _02068_ VPWR VGND _01080_ sg13g2_mux2_1
X_20442_ \atbs_core_0.spike_memory_0.n2359_o[1]\ VPWR VGND _02069_ sg13g2_buf_1
X_20443_ _02069_ \atbs_core_0.spike_memory_0.n2358_o[1]\ _02068_ VPWR VGND _01081_ sg13g2_mux2_1
X_20444_ \atbs_core_0.spike_memory_0.n2369_o[1]\ _02048_ _02068_ VPWR VGND _01082_ sg13g2_mux2_1
X_20445_ \atbs_core_0.spike_memory_0.n2369_o[2]\ _02049_ _02068_ VPWR VGND _01083_ sg13g2_mux2_1
X_20446_ \atbs_core_0.spike_memory_0.n2369_o[3]\ _02050_ _02068_ VPWR VGND _01084_ sg13g2_mux2_1
X_20447_ \atbs_core_0.spike_memory_0.n2369_o[4]\ _02051_ _02068_ VPWR VGND _01085_ sg13g2_mux2_1
X_20448_ \atbs_core_0.spike_memory_0.n2369_o[5]\ _02052_ _02068_ VPWR VGND _01086_ sg13g2_mux2_1
X_20449_ \atbs_core_0.spike_memory_0.n2369_o[6]\ _02053_ _02068_ VPWR VGND _01087_ sg13g2_mux2_1
X_20450_ \atbs_core_0.spike_memory_0.n2369_o[7]\ _02054_ _02068_ VPWR VGND _01088_ sg13g2_mux2_1
X_20451_ _02026_ VPWR VGND _02070_ sg13g2_buf_1
X_20452_ \atbs_core_0.spike_memory_0.n2369_o[8]\ _02055_ _02070_ VPWR VGND _01089_ sg13g2_mux2_1
X_20453_ \atbs_core_0.spike_memory_0.n2369_o[9]\ _02056_ _02070_ VPWR VGND _01090_ sg13g2_mux2_1
X_20454_ \atbs_core_0.spike_memory_0.n2369_o[10]\ _02059_ _02070_ VPWR VGND _01091_ sg13g2_mux2_1
X_20455_ \atbs_core_0.spike_memory_0.n2359_o[2]\ VPWR VGND _02071_ sg13g2_buf_1
X_20456_ _02071_ \atbs_core_0.spike_memory_0.n2358_o[2]\ _02070_ VPWR VGND _01092_ sg13g2_mux2_1
X_20457_ \atbs_core_0.spike_memory_0.n2369_o[11]\ _02060_ _02070_ VPWR VGND _01093_ sg13g2_mux2_1
X_20458_ \atbs_core_0.spike_memory_0.n2369_o[12]\ _02061_ _02070_ VPWR VGND _01094_ sg13g2_mux2_1
X_20459_ \atbs_core_0.spike_memory_0.n2369_o[13]\ _02062_ _02070_ VPWR VGND _01095_ sg13g2_mux2_1
X_20460_ \atbs_core_0.spike_memory_0.n2369_o[14]\ _02063_ _02070_ VPWR VGND _01096_ sg13g2_mux2_1
X_20461_ \atbs_core_0.spike_memory_0.n2369_o[15]\ _02064_ _02070_ VPWR VGND _01097_ sg13g2_mux2_1
X_20462_ \atbs_core_0.spike_memory_0.n2369_o[16]\ _02065_ _02070_ VPWR VGND _01098_ sg13g2_mux2_1
X_20463_ _02026_ VPWR VGND _02072_ sg13g2_buf_1
X_20464_ \atbs_core_0.spike_memory_0.n2369_o[17]\ _02066_ _02072_ VPWR VGND _01099_ sg13g2_mux2_1
X_20465_ \atbs_core_0.spike_memory_0.n2369_o[18]\ _02067_ _02072_ VPWR VGND _01100_ sg13g2_mux2_1
X_20466_ \atbs_core_0.spike_memory_0.n2370_o[0]\ \atbs_core_0.spike_memory_0.n2369_o[0]\ _02072_ VPWR VGND _01101_ sg13g2_mux2_1
X_20467_ \atbs_core_0.spike_memory_0.n2370_o[1]\ \atbs_core_0.spike_memory_0.n2369_o[1]\ _02072_ VPWR VGND _01102_ sg13g2_mux2_1
X_20468_ \atbs_core_0.spike_memory_0.n2359_o[3]\ VPWR VGND _02073_ sg13g2_buf_1
X_20469_ _02073_ \atbs_core_0.spike_memory_0.n2358_o[3]\ _02072_ VPWR VGND _01103_ sg13g2_mux2_1
X_20470_ \atbs_core_0.spike_memory_0.n2370_o[2]\ \atbs_core_0.spike_memory_0.n2369_o[2]\ _02072_ VPWR VGND _01104_ sg13g2_mux2_1
X_20471_ \atbs_core_0.spike_memory_0.n2370_o[3]\ \atbs_core_0.spike_memory_0.n2369_o[3]\ _02072_ VPWR VGND _01105_ sg13g2_mux2_1
X_20472_ \atbs_core_0.spike_memory_0.n2370_o[4]\ \atbs_core_0.spike_memory_0.n2369_o[4]\ _02072_ VPWR VGND _01106_ sg13g2_mux2_1
X_20473_ \atbs_core_0.spike_memory_0.n2370_o[5]\ \atbs_core_0.spike_memory_0.n2369_o[5]\ _02072_ VPWR VGND _01107_ sg13g2_mux2_1
X_20474_ \atbs_core_0.spike_memory_0.n2370_o[6]\ \atbs_core_0.spike_memory_0.n2369_o[6]\ _02072_ VPWR VGND _01108_ sg13g2_mux2_1
X_20475_ _12511_ VPWR VGND _02074_ sg13g2_buf_1
X_20476_ _02074_ VPWR VGND _02075_ sg13g2_buf_1
X_20477_ _02075_ VPWR VGND _02076_ sg13g2_buf_1
X_20478_ \atbs_core_0.spike_memory_0.n2370_o[7]\ \atbs_core_0.spike_memory_0.n2369_o[7]\ _02076_ VPWR VGND _01109_ sg13g2_mux2_1
X_20479_ \atbs_core_0.spike_memory_0.n2370_o[8]\ \atbs_core_0.spike_memory_0.n2369_o[8]\ _02076_ VPWR VGND _01110_ sg13g2_mux2_1
X_20480_ \atbs_core_0.spike_memory_0.n2370_o[9]\ \atbs_core_0.spike_memory_0.n2369_o[9]\ _02076_ VPWR VGND _01111_ sg13g2_mux2_1
X_20481_ \atbs_core_0.spike_memory_0.n2370_o[10]\ \atbs_core_0.spike_memory_0.n2369_o[10]\ _02076_ VPWR VGND _01112_ sg13g2_mux2_1
X_20482_ \atbs_core_0.spike_memory_0.n2370_o[11]\ \atbs_core_0.spike_memory_0.n2369_o[11]\ _02076_ VPWR VGND _01113_ sg13g2_mux2_1
X_20483_ \atbs_core_0.spike_memory_0.n2359_o[4]\ VPWR VGND _02077_ sg13g2_buf_1
X_20484_ _02077_ \atbs_core_0.spike_memory_0.n2358_o[4]\ _02076_ VPWR VGND _01114_ sg13g2_mux2_1
X_20485_ \atbs_core_0.spike_memory_0.n2370_o[12]\ \atbs_core_0.spike_memory_0.n2369_o[12]\ _02076_ VPWR VGND _01115_ sg13g2_mux2_1
X_20486_ \atbs_core_0.spike_memory_0.n2370_o[13]\ \atbs_core_0.spike_memory_0.n2369_o[13]\ _02076_ VPWR VGND _01116_ sg13g2_mux2_1
X_20487_ \atbs_core_0.spike_memory_0.n2370_o[14]\ \atbs_core_0.spike_memory_0.n2369_o[14]\ _02076_ VPWR VGND _01117_ sg13g2_mux2_1
X_20488_ \atbs_core_0.spike_memory_0.n2370_o[15]\ \atbs_core_0.spike_memory_0.n2369_o[15]\ _02076_ VPWR VGND _01118_ sg13g2_mux2_1
X_20489_ _02075_ VPWR VGND _02078_ sg13g2_buf_1
X_20490_ \atbs_core_0.spike_memory_0.n2370_o[16]\ \atbs_core_0.spike_memory_0.n2369_o[16]\ _02078_ VPWR VGND _01119_ sg13g2_mux2_1
X_20491_ \atbs_core_0.spike_memory_0.n2370_o[17]\ \atbs_core_0.spike_memory_0.n2369_o[17]\ _02078_ VPWR VGND _01120_ sg13g2_mux2_1
X_20492_ \atbs_core_0.spike_memory_0.n2370_o[18]\ \atbs_core_0.spike_memory_0.n2369_o[18]\ _02078_ VPWR VGND _01121_ sg13g2_mux2_1
X_20493_ \atbs_core_0.spike_memory_0.n2371_o[0]\ VPWR VGND _02079_ sg13g2_buf_1
X_20494_ _02079_ \atbs_core_0.spike_memory_0.n2370_o[0]\ _02078_ VPWR VGND _01122_ sg13g2_mux2_1
X_20495_ \atbs_core_0.spike_memory_0.n2371_o[1]\ VPWR VGND _02080_ sg13g2_buf_1
X_20496_ _02080_ \atbs_core_0.spike_memory_0.n2370_o[1]\ _02078_ VPWR VGND _01123_ sg13g2_mux2_1
X_20497_ \atbs_core_0.spike_memory_0.n2371_o[2]\ VPWR VGND _02081_ sg13g2_buf_1
X_20498_ _02081_ \atbs_core_0.spike_memory_0.n2370_o[2]\ _02078_ VPWR VGND _01124_ sg13g2_mux2_1
X_20499_ \atbs_core_0.spike_memory_0.n2359_o[5]\ VPWR VGND _02082_ sg13g2_buf_1
X_20500_ _02082_ \atbs_core_0.spike_memory_0.n2358_o[5]\ _02078_ VPWR VGND _01125_ sg13g2_mux2_1
X_20501_ \atbs_core_0.spike_memory_0.n2371_o[3]\ VPWR VGND _02083_ sg13g2_buf_1
X_20502_ _02083_ \atbs_core_0.spike_memory_0.n2370_o[3]\ _02078_ VPWR VGND _01126_ sg13g2_mux2_1
X_20503_ \atbs_core_0.spike_memory_0.n2371_o[4]\ VPWR VGND _02084_ sg13g2_buf_1
X_20504_ _02084_ \atbs_core_0.spike_memory_0.n2370_o[4]\ _02078_ VPWR VGND _01127_ sg13g2_mux2_1
X_20505_ \atbs_core_0.spike_memory_0.n2371_o[5]\ VPWR VGND _02085_ sg13g2_buf_1
X_20506_ _02085_ \atbs_core_0.spike_memory_0.n2370_o[5]\ _02078_ VPWR VGND _01128_ sg13g2_mux2_1
X_20507_ \atbs_core_0.spike_memory_0.n2371_o[6]\ VPWR VGND _02086_ sg13g2_buf_1
X_20508_ _02075_ VPWR VGND _02087_ sg13g2_buf_1
X_20509_ _02086_ \atbs_core_0.spike_memory_0.n2370_o[6]\ _02087_ VPWR VGND _01129_ sg13g2_mux2_1
X_20510_ \atbs_core_0.spike_memory_0.n2371_o[7]\ VPWR VGND _02088_ sg13g2_buf_1
X_20511_ _02088_ \atbs_core_0.spike_memory_0.n2370_o[7]\ _02087_ VPWR VGND _01130_ sg13g2_mux2_1
X_20512_ \atbs_core_0.spike_memory_0.n2371_o[8]\ VPWR VGND _02089_ sg13g2_buf_1
X_20513_ _02089_ \atbs_core_0.spike_memory_0.n2370_o[8]\ _02087_ VPWR VGND _01131_ sg13g2_mux2_1
X_20514_ \atbs_core_0.spike_memory_0.n2371_o[9]\ VPWR VGND _02090_ sg13g2_buf_1
X_20515_ _02090_ \atbs_core_0.spike_memory_0.n2370_o[9]\ _02087_ VPWR VGND _01132_ sg13g2_mux2_1
X_20516_ \atbs_core_0.spike_memory_0.n2371_o[10]\ VPWR VGND _02091_ sg13g2_buf_1
X_20517_ _02091_ \atbs_core_0.spike_memory_0.n2370_o[10]\ _02087_ VPWR VGND _01133_ sg13g2_mux2_1
X_20518_ \atbs_core_0.spike_memory_0.n2371_o[11]\ VPWR VGND _02092_ sg13g2_buf_1
X_20519_ _02092_ \atbs_core_0.spike_memory_0.n2370_o[11]\ _02087_ VPWR VGND _01134_ sg13g2_mux2_1
X_20520_ \atbs_core_0.spike_memory_0.n2371_o[12]\ VPWR VGND _02093_ sg13g2_buf_1
X_20521_ _02093_ \atbs_core_0.spike_memory_0.n2370_o[12]\ _02087_ VPWR VGND _01135_ sg13g2_mux2_1
X_20522_ \atbs_core_0.spike_memory_0.n2359_o[6]\ VPWR VGND _02094_ sg13g2_buf_1
X_20523_ _02094_ \atbs_core_0.spike_memory_0.n2358_o[6]\ _02087_ VPWR VGND _01136_ sg13g2_mux2_1
X_20524_ \atbs_core_0.spike_memory_0.n2371_o[13]\ VPWR VGND _02095_ sg13g2_buf_1
X_20525_ _02095_ \atbs_core_0.spike_memory_0.n2370_o[13]\ _02087_ VPWR VGND _01137_ sg13g2_mux2_1
X_20526_ \atbs_core_0.spike_memory_0.n2371_o[14]\ VPWR VGND _02096_ sg13g2_buf_1
X_20527_ _02096_ \atbs_core_0.spike_memory_0.n2370_o[14]\ _02087_ VPWR VGND _01138_ sg13g2_mux2_1
X_20528_ \atbs_core_0.spike_memory_0.n2371_o[15]\ VPWR VGND _02097_ sg13g2_buf_1
X_20529_ _02075_ VPWR VGND _02098_ sg13g2_buf_1
X_20530_ _02097_ \atbs_core_0.spike_memory_0.n2370_o[15]\ _02098_ VPWR VGND _01139_ sg13g2_mux2_1
X_20531_ \atbs_core_0.spike_memory_0.n2371_o[16]\ VPWR VGND _02099_ sg13g2_buf_1
X_20532_ _02099_ \atbs_core_0.spike_memory_0.n2370_o[16]\ _02098_ VPWR VGND _01140_ sg13g2_mux2_1
X_20533_ \atbs_core_0.spike_memory_0.n2371_o[17]\ VPWR VGND _02100_ sg13g2_buf_1
X_20534_ _02100_ \atbs_core_0.spike_memory_0.n2370_o[17]\ _02098_ VPWR VGND _01141_ sg13g2_mux2_1
X_20535_ \atbs_core_0.spike_memory_0.n2371_o[18]\ VPWR VGND _02101_ sg13g2_buf_1
X_20536_ _02101_ \atbs_core_0.spike_memory_0.n2370_o[18]\ _02098_ VPWR VGND _01142_ sg13g2_mux2_1
X_20537_ \atbs_core_0.spike_memory_0.n2372_o[0]\ VPWR VGND _02102_ sg13g2_buf_1
X_20538_ _02102_ _02079_ _02098_ VPWR VGND _01143_ sg13g2_mux2_1
X_20539_ \atbs_core_0.spike_memory_0.n2372_o[1]\ VPWR VGND _02103_ sg13g2_buf_1
X_20540_ _02103_ _02080_ _02098_ VPWR VGND _01144_ sg13g2_mux2_1
X_20541_ \atbs_core_0.spike_memory_0.n2372_o[2]\ VPWR VGND _02104_ sg13g2_buf_1
X_20542_ _02104_ _02081_ _02098_ VPWR VGND _01145_ sg13g2_mux2_1
X_20543_ \atbs_core_0.spike_memory_0.n2372_o[3]\ VPWR VGND _02105_ sg13g2_buf_1
X_20544_ _02105_ _02083_ _02098_ VPWR VGND _01146_ sg13g2_mux2_1
X_20545_ \atbs_core_0.spike_memory_0.n2359_o[7]\ VPWR VGND _02106_ sg13g2_buf_1
X_20546_ _02106_ \atbs_core_0.spike_memory_0.n2358_o[7]\ _02098_ VPWR VGND _01147_ sg13g2_mux2_1
X_20547_ \atbs_core_0.spike_memory_0.n2372_o[4]\ VPWR VGND _02107_ sg13g2_buf_1
X_20548_ _02107_ _02084_ _02098_ VPWR VGND _01148_ sg13g2_mux2_1
X_20549_ \atbs_core_0.spike_memory_0.n2372_o[5]\ VPWR VGND _02108_ sg13g2_buf_1
X_20550_ _02075_ VPWR VGND _02109_ sg13g2_buf_1
X_20551_ _02108_ _02085_ _02109_ VPWR VGND _01149_ sg13g2_mux2_1
X_20552_ \atbs_core_0.spike_memory_0.n2372_o[6]\ VPWR VGND _02110_ sg13g2_buf_1
X_20553_ _02110_ _02086_ _02109_ VPWR VGND _01150_ sg13g2_mux2_1
X_20554_ \atbs_core_0.spike_memory_0.n2372_o[7]\ VPWR VGND _02111_ sg13g2_buf_1
X_20555_ _02111_ _02088_ _02109_ VPWR VGND _01151_ sg13g2_mux2_1
X_20556_ \atbs_core_0.spike_memory_0.n2372_o[8]\ VPWR VGND _02112_ sg13g2_buf_1
X_20557_ _02112_ _02089_ _02109_ VPWR VGND _01152_ sg13g2_mux2_1
X_20558_ \atbs_core_0.spike_memory_0.n2372_o[9]\ VPWR VGND _02113_ sg13g2_buf_1
X_20559_ _02113_ _02090_ _02109_ VPWR VGND _01153_ sg13g2_mux2_1
X_20560_ \atbs_core_0.spike_memory_0.n2372_o[10]\ VPWR VGND _02114_ sg13g2_buf_1
X_20561_ _02114_ _02091_ _02109_ VPWR VGND _01154_ sg13g2_mux2_1
X_20562_ \atbs_core_0.spike_memory_0.n2372_o[11]\ VPWR VGND _02115_ sg13g2_buf_1
X_20563_ _02115_ _02092_ _02109_ VPWR VGND _01155_ sg13g2_mux2_1
X_20564_ \atbs_core_0.spike_memory_0.n2372_o[12]\ VPWR VGND _02116_ sg13g2_buf_1
X_20565_ _02116_ _02093_ _02109_ VPWR VGND _01156_ sg13g2_mux2_1
X_20566_ \atbs_core_0.spike_memory_0.n2372_o[13]\ VPWR VGND _02117_ sg13g2_buf_1
X_20567_ _02117_ _02095_ _02109_ VPWR VGND _01157_ sg13g2_mux2_1
X_20568_ \atbs_core_0.spike_memory_0.n2359_o[8]\ VPWR VGND _02118_ sg13g2_buf_1
X_20569_ _02118_ \atbs_core_0.spike_memory_0.n2358_o[8]\ _02109_ VPWR VGND _01158_ sg13g2_mux2_1
X_20570_ \atbs_core_0.spike_memory_0.n2372_o[14]\ VPWR VGND _02119_ sg13g2_buf_1
X_20571_ _02075_ VPWR VGND _02120_ sg13g2_buf_1
X_20572_ _02119_ _02096_ _02120_ VPWR VGND _01159_ sg13g2_mux2_1
X_20573_ \atbs_core_0.spike_memory_0.n2372_o[15]\ VPWR VGND _02121_ sg13g2_buf_1
X_20574_ _02121_ _02097_ _02120_ VPWR VGND _01160_ sg13g2_mux2_1
X_20575_ \atbs_core_0.spike_memory_0.n2372_o[16]\ VPWR VGND _02122_ sg13g2_buf_1
X_20576_ _02122_ _02099_ _02120_ VPWR VGND _01161_ sg13g2_mux2_1
X_20577_ \atbs_core_0.spike_memory_0.n2372_o[17]\ VPWR VGND _02123_ sg13g2_buf_1
X_20578_ _02123_ _02100_ _02120_ VPWR VGND _01162_ sg13g2_mux2_1
X_20579_ \atbs_core_0.spike_memory_0.n2372_o[18]\ VPWR VGND _02124_ sg13g2_buf_1
X_20580_ _02124_ _02101_ _02120_ VPWR VGND _01163_ sg13g2_mux2_1
X_20581_ \atbs_core_0.spike_memory_0.n2373_o[0]\ _02102_ _02120_ VPWR VGND _01164_ sg13g2_mux2_1
X_20582_ \atbs_core_0.spike_memory_0.n2373_o[1]\ _02103_ _02120_ VPWR VGND _01165_ sg13g2_mux2_1
X_20583_ \atbs_core_0.spike_memory_0.n2373_o[2]\ _02104_ _02120_ VPWR VGND _01166_ sg13g2_mux2_1
X_20584_ \atbs_core_0.spike_memory_0.n2373_o[3]\ _02105_ _02120_ VPWR VGND _01167_ sg13g2_mux2_1
X_20585_ \atbs_core_0.spike_memory_0.n2373_o[4]\ _02107_ _02120_ VPWR VGND _01168_ sg13g2_mux2_1
X_20586_ \atbs_core_0.spike_memory_0.n2359_o[9]\ VPWR VGND _02125_ sg13g2_buf_1
X_20587_ _02075_ VPWR VGND _02126_ sg13g2_buf_1
X_20588_ _02125_ \atbs_core_0.spike_memory_0.n2358_o[9]\ _02126_ VPWR VGND _01169_ sg13g2_mux2_1
X_20589_ \atbs_core_0.spike_memory_0.n2373_o[5]\ _02108_ _02126_ VPWR VGND _01170_ sg13g2_mux2_1
X_20590_ \atbs_core_0.spike_memory_0.n2373_o[6]\ _02110_ _02126_ VPWR VGND _01171_ sg13g2_mux2_1
X_20591_ \atbs_core_0.spike_memory_0.n2373_o[7]\ _02111_ _02126_ VPWR VGND _01172_ sg13g2_mux2_1
X_20592_ \atbs_core_0.spike_memory_0.n2373_o[8]\ _02112_ _02126_ VPWR VGND _01173_ sg13g2_mux2_1
X_20593_ \atbs_core_0.spike_memory_0.n2373_o[9]\ _02113_ _02126_ VPWR VGND _01174_ sg13g2_mux2_1
X_20594_ \atbs_core_0.spike_memory_0.n2373_o[10]\ _02114_ _02126_ VPWR VGND _01175_ sg13g2_mux2_1
X_20595_ \atbs_core_0.spike_memory_0.n2373_o[11]\ _02115_ _02126_ VPWR VGND _01176_ sg13g2_mux2_1
X_20596_ \atbs_core_0.spike_memory_0.n2373_o[12]\ _02116_ _02126_ VPWR VGND _01177_ sg13g2_mux2_1
X_20597_ \atbs_core_0.spike_memory_0.n2373_o[13]\ _02117_ _02126_ VPWR VGND _01178_ sg13g2_mux2_1
X_20598_ _02074_ VPWR VGND _02127_ sg13g2_buf_1
X_20599_ _02127_ VPWR VGND _02128_ sg13g2_buf_1
X_20600_ \atbs_core_0.spike_memory_0.n2373_o[14]\ _02119_ _02128_ VPWR VGND _01179_ sg13g2_mux2_1
X_20601_ \atbs_core_0.spike_memory_0.n2359_o[10]\ VPWR VGND _02129_ sg13g2_buf_1
X_20602_ _02129_ \atbs_core_0.spike_memory_0.n2358_o[10]\ _02128_ VPWR VGND _01180_ sg13g2_mux2_1
X_20603_ \atbs_core_0.spike_memory_0.n2358_o[2]\ \atbs_core_0.spike_memory_0.a_data[2]\ _02128_ VPWR VGND _01181_ sg13g2_mux2_1
X_20604_ \atbs_core_0.spike_memory_0.n2373_o[15]\ _02121_ _02128_ VPWR VGND _01182_ sg13g2_mux2_1
X_20605_ \atbs_core_0.spike_memory_0.n2373_o[16]\ _02122_ _02128_ VPWR VGND _01183_ sg13g2_mux2_1
X_20606_ \atbs_core_0.spike_memory_0.n2373_o[17]\ _02123_ _02128_ VPWR VGND _01184_ sg13g2_mux2_1
X_20607_ \atbs_core_0.spike_memory_0.n2373_o[18]\ _02124_ _02128_ VPWR VGND _01185_ sg13g2_mux2_1
X_20608_ \atbs_core_0.spike_memory_0.n2374_o[0]\ \atbs_core_0.spike_memory_0.n2373_o[0]\ _02128_ VPWR VGND _01186_ sg13g2_mux2_1
X_20609_ \atbs_core_0.spike_memory_0.n2374_o[1]\ \atbs_core_0.spike_memory_0.n2373_o[1]\ _02128_ VPWR VGND _01187_ sg13g2_mux2_1
X_20610_ \atbs_core_0.spike_memory_0.n2374_o[2]\ \atbs_core_0.spike_memory_0.n2373_o[2]\ _02128_ VPWR VGND _01188_ sg13g2_mux2_1
X_20611_ _02127_ VPWR VGND _02130_ sg13g2_buf_1
X_20612_ \atbs_core_0.spike_memory_0.n2374_o[3]\ \atbs_core_0.spike_memory_0.n2373_o[3]\ _02130_ VPWR VGND _01189_ sg13g2_mux2_1
X_20613_ \atbs_core_0.spike_memory_0.n2374_o[4]\ \atbs_core_0.spike_memory_0.n2373_o[4]\ _02130_ VPWR VGND _01190_ sg13g2_mux2_1
X_20614_ \atbs_core_0.spike_memory_0.n2374_o[5]\ \atbs_core_0.spike_memory_0.n2373_o[5]\ _02130_ VPWR VGND _01191_ sg13g2_mux2_1
X_20615_ \atbs_core_0.spike_memory_0.n2359_o[11]\ VPWR VGND _02131_ sg13g2_buf_1
X_20616_ _02131_ \atbs_core_0.spike_memory_0.n2358_o[11]\ _02130_ VPWR VGND _01192_ sg13g2_mux2_1
X_20617_ \atbs_core_0.spike_memory_0.n2374_o[6]\ \atbs_core_0.spike_memory_0.n2373_o[6]\ _02130_ VPWR VGND _01193_ sg13g2_mux2_1
X_20618_ \atbs_core_0.spike_memory_0.n2374_o[7]\ \atbs_core_0.spike_memory_0.n2373_o[7]\ _02130_ VPWR VGND _01194_ sg13g2_mux2_1
X_20619_ \atbs_core_0.spike_memory_0.n2374_o[8]\ \atbs_core_0.spike_memory_0.n2373_o[8]\ _02130_ VPWR VGND _01195_ sg13g2_mux2_1
X_20620_ \atbs_core_0.spike_memory_0.n2374_o[9]\ \atbs_core_0.spike_memory_0.n2373_o[9]\ _02130_ VPWR VGND _01196_ sg13g2_mux2_1
X_20621_ \atbs_core_0.spike_memory_0.n2374_o[10]\ \atbs_core_0.spike_memory_0.n2373_o[10]\ _02130_ VPWR VGND _01197_ sg13g2_mux2_1
X_20622_ \atbs_core_0.spike_memory_0.n2374_o[11]\ \atbs_core_0.spike_memory_0.n2373_o[11]\ _02130_ VPWR VGND _01198_ sg13g2_mux2_1
X_20623_ _02127_ VPWR VGND _02132_ sg13g2_buf_1
X_20624_ \atbs_core_0.spike_memory_0.n2374_o[12]\ \atbs_core_0.spike_memory_0.n2373_o[12]\ _02132_ VPWR VGND _01199_ sg13g2_mux2_1
X_20625_ \atbs_core_0.spike_memory_0.n2374_o[13]\ \atbs_core_0.spike_memory_0.n2373_o[13]\ _02132_ VPWR VGND _01200_ sg13g2_mux2_1
X_20626_ \atbs_core_0.spike_memory_0.n2374_o[14]\ \atbs_core_0.spike_memory_0.n2373_o[14]\ _02132_ VPWR VGND _01201_ sg13g2_mux2_1
X_20627_ \atbs_core_0.spike_memory_0.n2374_o[15]\ \atbs_core_0.spike_memory_0.n2373_o[15]\ _02132_ VPWR VGND _01202_ sg13g2_mux2_1
X_20628_ \atbs_core_0.spike_memory_0.n2359_o[12]\ VPWR VGND _02133_ sg13g2_buf_1
X_20629_ _02133_ \atbs_core_0.spike_memory_0.n2358_o[12]\ _02132_ VPWR VGND _01203_ sg13g2_mux2_1
X_20630_ \atbs_core_0.spike_memory_0.n2374_o[16]\ \atbs_core_0.spike_memory_0.n2373_o[16]\ _02132_ VPWR VGND _01204_ sg13g2_mux2_1
X_20631_ \atbs_core_0.spike_memory_0.n2374_o[17]\ \atbs_core_0.spike_memory_0.n2373_o[17]\ _02132_ VPWR VGND _01205_ sg13g2_mux2_1
X_20632_ \atbs_core_0.spike_memory_0.n2374_o[18]\ \atbs_core_0.spike_memory_0.n2373_o[18]\ _02132_ VPWR VGND _01206_ sg13g2_mux2_1
X_20633_ \atbs_core_0.spike_memory_0.n2375_o[0]\ VPWR VGND _02134_ sg13g2_buf_1
X_20634_ _02134_ \atbs_core_0.spike_memory_0.n2374_o[0]\ _02132_ VPWR VGND _01207_ sg13g2_mux2_1
X_20635_ \atbs_core_0.spike_memory_0.n2375_o[1]\ VPWR VGND _02135_ sg13g2_buf_1
X_20636_ _02135_ \atbs_core_0.spike_memory_0.n2374_o[1]\ _02132_ VPWR VGND _01208_ sg13g2_mux2_1
X_20637_ \atbs_core_0.spike_memory_0.n2375_o[2]\ VPWR VGND _02136_ sg13g2_buf_1
X_20638_ _02127_ VPWR VGND _02137_ sg13g2_buf_1
X_20639_ _02136_ \atbs_core_0.spike_memory_0.n2374_o[2]\ _02137_ VPWR VGND _01209_ sg13g2_mux2_1
X_20640_ \atbs_core_0.spike_memory_0.n2375_o[3]\ VPWR VGND _02138_ sg13g2_buf_1
X_20641_ _02138_ \atbs_core_0.spike_memory_0.n2374_o[3]\ _02137_ VPWR VGND _01210_ sg13g2_mux2_1
X_20642_ \atbs_core_0.spike_memory_0.n2375_o[4]\ VPWR VGND _02139_ sg13g2_buf_1
X_20643_ _02139_ \atbs_core_0.spike_memory_0.n2374_o[4]\ _02137_ VPWR VGND _01211_ sg13g2_mux2_1
X_20644_ \atbs_core_0.spike_memory_0.n2375_o[5]\ VPWR VGND _02140_ sg13g2_buf_1
X_20645_ _02140_ \atbs_core_0.spike_memory_0.n2374_o[5]\ _02137_ VPWR VGND _01212_ sg13g2_mux2_1
X_20646_ \atbs_core_0.spike_memory_0.n2375_o[6]\ VPWR VGND _02141_ sg13g2_buf_1
X_20647_ _02141_ \atbs_core_0.spike_memory_0.n2374_o[6]\ _02137_ VPWR VGND _01213_ sg13g2_mux2_1
X_20648_ \atbs_core_0.spike_memory_0.n2359_o[13]\ VPWR VGND _02142_ sg13g2_buf_1
X_20649_ _02142_ \atbs_core_0.spike_memory_0.n2358_o[13]\ _02137_ VPWR VGND _01214_ sg13g2_mux2_1
X_20650_ \atbs_core_0.spike_memory_0.n2375_o[7]\ VPWR VGND _02143_ sg13g2_buf_1
X_20651_ _02143_ \atbs_core_0.spike_memory_0.n2374_o[7]\ _02137_ VPWR VGND _01215_ sg13g2_mux2_1
X_20652_ \atbs_core_0.spike_memory_0.n2375_o[8]\ VPWR VGND _02144_ sg13g2_buf_1
X_20653_ _02144_ \atbs_core_0.spike_memory_0.n2374_o[8]\ _02137_ VPWR VGND _01216_ sg13g2_mux2_1
X_20654_ \atbs_core_0.spike_memory_0.n2375_o[9]\ VPWR VGND _02145_ sg13g2_buf_1
X_20655_ _02145_ \atbs_core_0.spike_memory_0.n2374_o[9]\ _02137_ VPWR VGND _01217_ sg13g2_mux2_1
X_20656_ \atbs_core_0.spike_memory_0.n2375_o[10]\ VPWR VGND _02146_ sg13g2_buf_1
X_20657_ _02146_ \atbs_core_0.spike_memory_0.n2374_o[10]\ _02137_ VPWR VGND _01218_ sg13g2_mux2_1
X_20658_ \atbs_core_0.spike_memory_0.n2375_o[11]\ VPWR VGND _02147_ sg13g2_buf_1
X_20659_ _02127_ VPWR VGND _02148_ sg13g2_buf_1
X_20660_ _02147_ \atbs_core_0.spike_memory_0.n2374_o[11]\ _02148_ VPWR VGND _01219_ sg13g2_mux2_1
X_20661_ \atbs_core_0.spike_memory_0.n2375_o[12]\ VPWR VGND _02149_ sg13g2_buf_1
X_20662_ _02149_ \atbs_core_0.spike_memory_0.n2374_o[12]\ _02148_ VPWR VGND _01220_ sg13g2_mux2_1
X_20663_ \atbs_core_0.spike_memory_0.n2375_o[13]\ VPWR VGND _02150_ sg13g2_buf_1
X_20664_ _02150_ \atbs_core_0.spike_memory_0.n2374_o[13]\ _02148_ VPWR VGND _01221_ sg13g2_mux2_1
X_20665_ \atbs_core_0.spike_memory_0.n2375_o[14]\ VPWR VGND _02151_ sg13g2_buf_1
X_20666_ _02151_ \atbs_core_0.spike_memory_0.n2374_o[14]\ _02148_ VPWR VGND _01222_ sg13g2_mux2_1
X_20667_ \atbs_core_0.spike_memory_0.n2375_o[15]\ VPWR VGND _02152_ sg13g2_buf_1
X_20668_ _02152_ \atbs_core_0.spike_memory_0.n2374_o[15]\ _02148_ VPWR VGND _01223_ sg13g2_mux2_1
X_20669_ \atbs_core_0.spike_memory_0.n2375_o[16]\ VPWR VGND _02153_ sg13g2_buf_1
X_20670_ _02153_ \atbs_core_0.spike_memory_0.n2374_o[16]\ _02148_ VPWR VGND _01224_ sg13g2_mux2_1
X_20671_ \atbs_core_0.spike_memory_0.n2359_o[14]\ VPWR VGND _02154_ sg13g2_buf_1
X_20672_ _02154_ \atbs_core_0.spike_memory_0.n2358_o[14]\ _02148_ VPWR VGND _01225_ sg13g2_mux2_1
X_20673_ \atbs_core_0.spike_memory_0.n2375_o[17]\ VPWR VGND _02155_ sg13g2_buf_1
X_20674_ _02155_ \atbs_core_0.spike_memory_0.n2374_o[17]\ _02148_ VPWR VGND _01226_ sg13g2_mux2_1
X_20675_ \atbs_core_0.spike_memory_0.n2375_o[18]\ VPWR VGND _02156_ sg13g2_buf_1
X_20676_ _02156_ \atbs_core_0.spike_memory_0.n2374_o[18]\ _02148_ VPWR VGND _01227_ sg13g2_mux2_1
X_20677_ \atbs_core_0.spike_memory_0.n2376_o[0]\ VPWR VGND _02157_ sg13g2_buf_1
X_20678_ _02157_ _02134_ _02148_ VPWR VGND _01228_ sg13g2_mux2_1
X_20679_ \atbs_core_0.spike_memory_0.n2376_o[1]\ VPWR VGND _02158_ sg13g2_buf_1
X_20680_ _02127_ VPWR VGND _02159_ sg13g2_buf_1
X_20681_ _02158_ _02135_ _02159_ VPWR VGND _01229_ sg13g2_mux2_1
X_20682_ \atbs_core_0.spike_memory_0.n2376_o[2]\ VPWR VGND _02160_ sg13g2_buf_1
X_20683_ _02160_ _02136_ _02159_ VPWR VGND _01230_ sg13g2_mux2_1
X_20684_ \atbs_core_0.spike_memory_0.n2376_o[3]\ VPWR VGND _02161_ sg13g2_buf_1
X_20685_ _02161_ _02138_ _02159_ VPWR VGND _01231_ sg13g2_mux2_1
X_20686_ \atbs_core_0.spike_memory_0.n2376_o[4]\ VPWR VGND _02162_ sg13g2_buf_1
X_20687_ _02162_ _02139_ _02159_ VPWR VGND _01232_ sg13g2_mux2_1
X_20688_ \atbs_core_0.spike_memory_0.n2376_o[5]\ VPWR VGND _02163_ sg13g2_buf_1
X_20689_ _02163_ _02140_ _02159_ VPWR VGND _01233_ sg13g2_mux2_1
X_20690_ \atbs_core_0.spike_memory_0.n2376_o[6]\ VPWR VGND _02164_ sg13g2_buf_1
X_20691_ _02164_ _02141_ _02159_ VPWR VGND _01234_ sg13g2_mux2_1
X_20692_ \atbs_core_0.spike_memory_0.n2376_o[7]\ VPWR VGND _02165_ sg13g2_buf_1
X_20693_ _02165_ _02143_ _02159_ VPWR VGND _01235_ sg13g2_mux2_1
X_20694_ \atbs_core_0.spike_memory_0.n2359_o[15]\ VPWR VGND _02166_ sg13g2_buf_1
X_20695_ _02166_ \atbs_core_0.spike_memory_0.n2358_o[15]\ _02159_ VPWR VGND _01236_ sg13g2_mux2_1
X_20696_ \atbs_core_0.spike_memory_0.n2376_o[8]\ VPWR VGND _02167_ sg13g2_buf_1
X_20697_ _02167_ _02144_ _02159_ VPWR VGND _01237_ sg13g2_mux2_1
X_20698_ \atbs_core_0.spike_memory_0.n2376_o[9]\ VPWR VGND _02168_ sg13g2_buf_1
X_20699_ _02168_ _02145_ _02159_ VPWR VGND _01238_ sg13g2_mux2_1
X_20700_ \atbs_core_0.spike_memory_0.n2376_o[10]\ VPWR VGND _02169_ sg13g2_buf_1
X_20701_ _02127_ VPWR VGND _02170_ sg13g2_buf_1
X_20702_ _02169_ _02146_ _02170_ VPWR VGND _01239_ sg13g2_mux2_1
X_20703_ \atbs_core_0.spike_memory_0.n2376_o[11]\ VPWR VGND _02171_ sg13g2_buf_1
X_20704_ _02171_ _02147_ _02170_ VPWR VGND _01240_ sg13g2_mux2_1
X_20705_ \atbs_core_0.spike_memory_0.n2376_o[12]\ VPWR VGND _02172_ sg13g2_buf_1
X_20706_ _02172_ _02149_ _02170_ VPWR VGND _01241_ sg13g2_mux2_1
X_20707_ \atbs_core_0.spike_memory_0.n2376_o[13]\ VPWR VGND _02173_ sg13g2_buf_1
X_20708_ _02173_ _02150_ _02170_ VPWR VGND _01242_ sg13g2_mux2_1
X_20709_ \atbs_core_0.spike_memory_0.n2376_o[14]\ VPWR VGND _02174_ sg13g2_buf_1
X_20710_ _02174_ _02151_ _02170_ VPWR VGND _01243_ sg13g2_mux2_1
X_20711_ \atbs_core_0.spike_memory_0.n2376_o[15]\ VPWR VGND _02175_ sg13g2_buf_1
X_20712_ _02175_ _02152_ _02170_ VPWR VGND _01244_ sg13g2_mux2_1
X_20713_ \atbs_core_0.spike_memory_0.n2376_o[16]\ VPWR VGND _02176_ sg13g2_buf_1
X_20714_ _02176_ _02153_ _02170_ VPWR VGND _01245_ sg13g2_mux2_1
X_20715_ \atbs_core_0.spike_memory_0.n2376_o[17]\ VPWR VGND _02177_ sg13g2_buf_1
X_20716_ _02177_ _02155_ _02170_ VPWR VGND _01246_ sg13g2_mux2_1
X_20717_ \atbs_core_0.spike_memory_0.n2359_o[16]\ VPWR VGND _02178_ sg13g2_buf_1
X_20718_ _02178_ \atbs_core_0.spike_memory_0.n2358_o[16]\ _02170_ VPWR VGND _01247_ sg13g2_mux2_1
X_20719_ \atbs_core_0.spike_memory_0.n2376_o[18]\ VPWR VGND _02179_ sg13g2_buf_1
X_20720_ _02179_ _02156_ _02170_ VPWR VGND _01248_ sg13g2_mux2_1
X_20721_ \atbs_core_0.spike_memory_0.n2377_o[0]\ VPWR VGND _02180_ sg13g2_inv_1
X_20722_ _12513_ VPWR VGND _02181_ sg13g2_buf_1
X_20723_ _12512_ VPWR VGND _02182_ sg13g2_buf_1
X_20724_ _02157_ _02182_ VPWR VGND _02183_ sg13g2_nand2_1
X_20725_ _02180_ _02181_ _02183_ VPWR VGND _01249_ sg13g2_o21ai_1
X_20726_ \atbs_core_0.spike_memory_0.n2377_o[1]\ VPWR VGND _02184_ sg13g2_inv_1
X_20727_ _02158_ _02182_ VPWR VGND _02185_ sg13g2_nand2_1
X_20728_ _02184_ _02181_ _02185_ VPWR VGND _01250_ sg13g2_o21ai_1
X_20729_ \atbs_core_0.spike_memory_0.n2377_o[2]\ VPWR VGND _02186_ sg13g2_inv_1
X_20730_ _02160_ _02182_ VPWR VGND _02187_ sg13g2_nand2_1
X_20731_ _02186_ _02181_ _02187_ VPWR VGND _01251_ sg13g2_o21ai_1
X_20732_ \atbs_core_0.spike_memory_0.n2377_o[3]\ VPWR VGND _02188_ sg13g2_inv_1
X_20733_ _02161_ _02182_ VPWR VGND _02189_ sg13g2_nand2_1
X_20734_ _02188_ _02181_ _02189_ VPWR VGND _01252_ sg13g2_o21ai_1
X_20735_ \atbs_core_0.spike_memory_0.n2377_o[4]\ VPWR VGND _02190_ sg13g2_inv_1
X_20736_ _12511_ VPWR VGND _02191_ sg13g2_buf_1
X_20737_ _02191_ VPWR VGND _02192_ sg13g2_buf_1
X_20738_ _02162_ _02192_ VPWR VGND _02193_ sg13g2_nand2_1
X_20739_ _02190_ _02181_ _02193_ VPWR VGND _01253_ sg13g2_o21ai_1
X_20740_ \atbs_core_0.spike_memory_0.n2377_o[5]\ VPWR VGND _02194_ sg13g2_inv_1
X_20741_ _02163_ _02192_ VPWR VGND _02195_ sg13g2_nand2_1
X_20742_ _02194_ _02181_ _02195_ VPWR VGND _01254_ sg13g2_o21ai_1
X_20743_ \atbs_core_0.spike_memory_0.n2377_o[6]\ VPWR VGND _02196_ sg13g2_inv_1
X_20744_ _02164_ _02192_ VPWR VGND _02197_ sg13g2_nand2_1
X_20745_ _02196_ _02181_ _02197_ VPWR VGND _01255_ sg13g2_o21ai_1
X_20746_ \atbs_core_0.spike_memory_0.n2377_o[7]\ VPWR VGND _02198_ sg13g2_inv_1
X_20747_ _02165_ _02192_ VPWR VGND _02199_ sg13g2_nand2_1
X_20748_ _02198_ _02181_ _02199_ VPWR VGND _01256_ sg13g2_o21ai_1
X_20749_ \atbs_core_0.spike_memory_0.n2377_o[8]\ VPWR VGND _02200_ sg13g2_inv_1
X_20750_ _02167_ _02192_ VPWR VGND _02201_ sg13g2_nand2_1
X_20751_ _02200_ _02181_ _02201_ VPWR VGND _01257_ sg13g2_o21ai_1
X_20752_ \atbs_core_0.spike_memory_0.n2359_o[17]\ VPWR VGND _02202_ sg13g2_buf_1
X_20753_ _02074_ VPWR VGND _02203_ sg13g2_buf_1
X_20754_ _02203_ VPWR VGND _02204_ sg13g2_buf_1
X_20755_ _02202_ \atbs_core_0.spike_memory_0.n2358_o[17]\ _02204_ VPWR VGND _01258_ sg13g2_mux2_1
X_20756_ \atbs_core_0.spike_memory_0.n2377_o[9]\ VPWR VGND _02205_ sg13g2_inv_1
X_20757_ _02168_ _02192_ VPWR VGND _02206_ sg13g2_nand2_1
X_20758_ _02205_ _02181_ _02206_ VPWR VGND _01259_ sg13g2_o21ai_1
X_20759_ \atbs_core_0.spike_memory_0.n2377_o[10]\ VPWR VGND _02207_ sg13g2_inv_1
X_20760_ _12513_ VPWR VGND _02208_ sg13g2_buf_1
X_20761_ _02169_ _02192_ VPWR VGND _02209_ sg13g2_nand2_1
X_20762_ _02207_ _02208_ _02209_ VPWR VGND _01260_ sg13g2_o21ai_1
X_20763_ \atbs_core_0.spike_memory_0.n2377_o[11]\ VPWR VGND _02210_ sg13g2_inv_1
X_20764_ _02171_ _02192_ VPWR VGND _02211_ sg13g2_nand2_1
X_20765_ _02210_ _02208_ _02211_ VPWR VGND _01261_ sg13g2_o21ai_1
X_20766_ \atbs_core_0.spike_memory_0.n2377_o[12]\ VPWR VGND _02212_ sg13g2_inv_1
X_20767_ _02172_ _02192_ VPWR VGND _02213_ sg13g2_nand2_1
X_20768_ _02212_ _02208_ _02213_ VPWR VGND _01262_ sg13g2_o21ai_1
X_20769_ \atbs_core_0.spike_memory_0.n2377_o[13]\ VPWR VGND _02214_ sg13g2_inv_1
X_20770_ _02173_ _02192_ VPWR VGND _02215_ sg13g2_nand2_1
X_20771_ _02214_ _02208_ _02215_ VPWR VGND _01263_ sg13g2_o21ai_1
X_20772_ \atbs_core_0.spike_memory_0.n2377_o[14]\ VPWR VGND _02216_ sg13g2_inv_1
X_20773_ _02191_ VPWR VGND _02217_ sg13g2_buf_1
X_20774_ _02174_ _02217_ VPWR VGND _02218_ sg13g2_nand2_1
X_20775_ _02216_ _02208_ _02218_ VPWR VGND _01264_ sg13g2_o21ai_1
X_20776_ \atbs_core_0.spike_memory_0.n2377_o[15]\ VPWR VGND _02219_ sg13g2_inv_1
X_20777_ _02175_ _02217_ VPWR VGND _02220_ sg13g2_nand2_1
X_20778_ _02219_ _02208_ _02220_ VPWR VGND _01265_ sg13g2_o21ai_1
X_20779_ \atbs_core_0.spike_memory_0.n2377_o[16]\ VPWR VGND _02221_ sg13g2_inv_1
X_20780_ _02176_ _02217_ VPWR VGND _02222_ sg13g2_nand2_1
X_20781_ _02221_ _02208_ _02222_ VPWR VGND _01266_ sg13g2_o21ai_1
X_20782_ \atbs_core_0.spike_memory_0.n2377_o[17]\ VPWR VGND _02223_ sg13g2_inv_1
X_20783_ _02177_ _02217_ VPWR VGND _02224_ sg13g2_nand2_1
X_20784_ _02223_ _02208_ _02224_ VPWR VGND _01267_ sg13g2_o21ai_1
X_20785_ \atbs_core_0.spike_memory_0.n2377_o[18]\ VPWR VGND _02225_ sg13g2_inv_1
X_20786_ _02179_ _02217_ VPWR VGND _02226_ sg13g2_nand2_1
X_20787_ _02225_ _02208_ _02226_ VPWR VGND _01268_ sg13g2_o21ai_1
X_20788_ \atbs_core_0.spike_memory_0.n2359_o[18]\ VPWR VGND _02227_ sg13g2_buf_1
X_20789_ _02227_ \atbs_core_0.spike_memory_0.n2358_o[18]\ _02204_ VPWR VGND _01269_ sg13g2_mux2_1
X_20790_ \atbs_core_0.spike_memory_0.n2378_o[0]\ \atbs_core_0.spike_memory_0.n2377_o[0]\ _02204_ VPWR VGND _01270_ sg13g2_mux2_1
X_20791_ \atbs_core_0.spike_memory_0.n2378_o[1]\ \atbs_core_0.spike_memory_0.n2377_o[1]\ _02204_ VPWR VGND _01271_ sg13g2_mux2_1
X_20792_ \atbs_core_0.spike_memory_0.n2378_o[2]\ \atbs_core_0.spike_memory_0.n2377_o[2]\ _02204_ VPWR VGND _01272_ sg13g2_mux2_1
X_20793_ \atbs_core_0.spike_memory_0.n2378_o[3]\ \atbs_core_0.spike_memory_0.n2377_o[3]\ _02204_ VPWR VGND _01273_ sg13g2_mux2_1
X_20794_ \atbs_core_0.spike_memory_0.n2378_o[4]\ \atbs_core_0.spike_memory_0.n2377_o[4]\ _02204_ VPWR VGND _01274_ sg13g2_mux2_1
X_20795_ \atbs_core_0.spike_memory_0.n2378_o[5]\ \atbs_core_0.spike_memory_0.n2377_o[5]\ _02204_ VPWR VGND _01275_ sg13g2_mux2_1
X_20796_ \atbs_core_0.spike_memory_0.n2378_o[6]\ \atbs_core_0.spike_memory_0.n2377_o[6]\ _02204_ VPWR VGND _01276_ sg13g2_mux2_1
X_20797_ \atbs_core_0.spike_memory_0.n2378_o[7]\ \atbs_core_0.spike_memory_0.n2377_o[7]\ _02204_ VPWR VGND _01277_ sg13g2_mux2_1
X_20798_ _02203_ VPWR VGND _02228_ sg13g2_buf_1
X_20799_ \atbs_core_0.spike_memory_0.n2378_o[8]\ \atbs_core_0.spike_memory_0.n2377_o[8]\ _02228_ VPWR VGND _01278_ sg13g2_mux2_1
X_20800_ \atbs_core_0.spike_memory_0.n2378_o[9]\ \atbs_core_0.spike_memory_0.n2377_o[9]\ _02228_ VPWR VGND _01279_ sg13g2_mux2_1
X_20801_ \atbs_core_0.spike_memory_0.n2360_o[0]\ VPWR VGND _02229_ sg13g2_buf_1
X_20802_ _02229_ _02057_ _02228_ VPWR VGND _01280_ sg13g2_mux2_1
X_20803_ \atbs_core_0.spike_memory_0.n2378_o[10]\ \atbs_core_0.spike_memory_0.n2377_o[10]\ _02228_ VPWR VGND _01281_ sg13g2_mux2_1
X_20804_ \atbs_core_0.spike_memory_0.n2378_o[11]\ \atbs_core_0.spike_memory_0.n2377_o[11]\ _02228_ VPWR VGND _01282_ sg13g2_mux2_1
X_20805_ \atbs_core_0.spike_memory_0.n2378_o[12]\ \atbs_core_0.spike_memory_0.n2377_o[12]\ _02228_ VPWR VGND _01283_ sg13g2_mux2_1
X_20806_ \atbs_core_0.spike_memory_0.n2378_o[13]\ \atbs_core_0.spike_memory_0.n2377_o[13]\ _02228_ VPWR VGND _01284_ sg13g2_mux2_1
X_20807_ \atbs_core_0.spike_memory_0.n2378_o[14]\ \atbs_core_0.spike_memory_0.n2377_o[14]\ _02228_ VPWR VGND _01285_ sg13g2_mux2_1
X_20808_ \atbs_core_0.spike_memory_0.n2378_o[15]\ \atbs_core_0.spike_memory_0.n2377_o[15]\ _02228_ VPWR VGND _01286_ sg13g2_mux2_1
X_20809_ \atbs_core_0.spike_memory_0.n2378_o[16]\ \atbs_core_0.spike_memory_0.n2377_o[16]\ _02228_ VPWR VGND _01287_ sg13g2_mux2_1
X_20810_ _02203_ VPWR VGND _02230_ sg13g2_buf_1
X_20811_ \atbs_core_0.spike_memory_0.n2378_o[17]\ \atbs_core_0.spike_memory_0.n2377_o[17]\ _02230_ VPWR VGND _01288_ sg13g2_mux2_1
X_20812_ \atbs_core_0.spike_memory_0.n2378_o[18]\ \atbs_core_0.spike_memory_0.n2377_o[18]\ _02230_ VPWR VGND _01289_ sg13g2_mux2_1
X_20813_ \atbs_core_0.spike_memory_0.n2379_o[0]\ VPWR VGND _02231_ sg13g2_buf_1
X_20814_ _02231_ \atbs_core_0.spike_memory_0.n2378_o[0]\ _02230_ VPWR VGND _01290_ sg13g2_mux2_1
X_20815_ \atbs_core_0.spike_memory_0.n2360_o[1]\ VPWR VGND _02232_ sg13g2_buf_1
X_20816_ _02232_ _02069_ _02230_ VPWR VGND _01291_ sg13g2_mux2_1
X_20817_ \atbs_core_0.spike_memory_0.n2358_o[3]\ \atbs_core_0.spike_memory_0.a_data[3]\ _02230_ VPWR VGND _01292_ sg13g2_mux2_1
X_20818_ \atbs_core_0.spike_memory_0.n2379_o[1]\ VPWR VGND _02233_ sg13g2_buf_1
X_20819_ _02233_ \atbs_core_0.spike_memory_0.n2378_o[1]\ _02230_ VPWR VGND _01293_ sg13g2_mux2_1
X_20820_ \atbs_core_0.spike_memory_0.n2379_o[2]\ VPWR VGND _02234_ sg13g2_buf_1
X_20821_ _02234_ \atbs_core_0.spike_memory_0.n2378_o[2]\ _02230_ VPWR VGND _01294_ sg13g2_mux2_1
X_20822_ \atbs_core_0.spike_memory_0.n2379_o[3]\ VPWR VGND _02235_ sg13g2_buf_1
X_20823_ _02235_ \atbs_core_0.spike_memory_0.n2378_o[3]\ _02230_ VPWR VGND _01295_ sg13g2_mux2_1
X_20824_ \atbs_core_0.spike_memory_0.n2379_o[4]\ VPWR VGND _02236_ sg13g2_buf_1
X_20825_ _02236_ \atbs_core_0.spike_memory_0.n2378_o[4]\ _02230_ VPWR VGND _01296_ sg13g2_mux2_1
X_20826_ \atbs_core_0.spike_memory_0.n2379_o[5]\ VPWR VGND _02237_ sg13g2_buf_1
X_20827_ _02237_ \atbs_core_0.spike_memory_0.n2378_o[5]\ _02230_ VPWR VGND _01297_ sg13g2_mux2_1
X_20828_ \atbs_core_0.spike_memory_0.n2379_o[6]\ VPWR VGND _02238_ sg13g2_buf_1
X_20829_ _02203_ VPWR VGND _02239_ sg13g2_buf_1
X_20830_ _02238_ \atbs_core_0.spike_memory_0.n2378_o[6]\ _02239_ VPWR VGND _01298_ sg13g2_mux2_1
X_20831_ \atbs_core_0.spike_memory_0.n2379_o[7]\ VPWR VGND _02240_ sg13g2_buf_1
X_20832_ _02240_ \atbs_core_0.spike_memory_0.n2378_o[7]\ _02239_ VPWR VGND _01299_ sg13g2_mux2_1
X_20833_ \atbs_core_0.spike_memory_0.n2379_o[8]\ VPWR VGND _02241_ sg13g2_buf_1
X_20834_ _02241_ \atbs_core_0.spike_memory_0.n2378_o[8]\ _02239_ VPWR VGND _01300_ sg13g2_mux2_1
X_20835_ \atbs_core_0.spike_memory_0.n2379_o[9]\ VPWR VGND _02242_ sg13g2_buf_1
X_20836_ _02242_ \atbs_core_0.spike_memory_0.n2378_o[9]\ _02239_ VPWR VGND _01301_ sg13g2_mux2_1
X_20837_ \atbs_core_0.spike_memory_0.n2379_o[10]\ VPWR VGND _02243_ sg13g2_buf_1
X_20838_ _02243_ \atbs_core_0.spike_memory_0.n2378_o[10]\ _02239_ VPWR VGND _01302_ sg13g2_mux2_1
X_20839_ \atbs_core_0.spike_memory_0.n2360_o[2]\ VPWR VGND _02244_ sg13g2_buf_1
X_20840_ _02244_ _02071_ _02239_ VPWR VGND _01303_ sg13g2_mux2_1
X_20841_ \atbs_core_0.spike_memory_0.n2379_o[11]\ VPWR VGND _02245_ sg13g2_buf_1
X_20842_ _02245_ \atbs_core_0.spike_memory_0.n2378_o[11]\ _02239_ VPWR VGND _01304_ sg13g2_mux2_1
X_20843_ \atbs_core_0.spike_memory_0.n2379_o[12]\ VPWR VGND _02246_ sg13g2_buf_1
X_20844_ _02246_ \atbs_core_0.spike_memory_0.n2378_o[12]\ _02239_ VPWR VGND _01305_ sg13g2_mux2_1
X_20845_ \atbs_core_0.spike_memory_0.n2379_o[13]\ VPWR VGND _02247_ sg13g2_buf_1
X_20846_ _02247_ \atbs_core_0.spike_memory_0.n2378_o[13]\ _02239_ VPWR VGND _01306_ sg13g2_mux2_1
X_20847_ \atbs_core_0.spike_memory_0.n2379_o[14]\ VPWR VGND _02248_ sg13g2_buf_1
X_20848_ _02248_ \atbs_core_0.spike_memory_0.n2378_o[14]\ _02239_ VPWR VGND _01307_ sg13g2_mux2_1
X_20849_ \atbs_core_0.spike_memory_0.n2379_o[15]\ VPWR VGND _02249_ sg13g2_buf_1
X_20850_ _02203_ VPWR VGND _02250_ sg13g2_buf_1
X_20851_ _02249_ \atbs_core_0.spike_memory_0.n2378_o[15]\ _02250_ VPWR VGND _01308_ sg13g2_mux2_1
X_20852_ \atbs_core_0.spike_memory_0.n2379_o[16]\ VPWR VGND _02251_ sg13g2_buf_1
X_20853_ _02251_ \atbs_core_0.spike_memory_0.n2378_o[16]\ _02250_ VPWR VGND _01309_ sg13g2_mux2_1
X_20854_ \atbs_core_0.spike_memory_0.n2379_o[17]\ VPWR VGND _02252_ sg13g2_buf_1
X_20855_ _02252_ \atbs_core_0.spike_memory_0.n2378_o[17]\ _02250_ VPWR VGND _01310_ sg13g2_mux2_1
X_20856_ \atbs_core_0.spike_memory_0.n2379_o[18]\ VPWR VGND _02253_ sg13g2_buf_1
X_20857_ _02253_ \atbs_core_0.spike_memory_0.n2378_o[18]\ _02250_ VPWR VGND _01311_ sg13g2_mux2_1
X_20858_ \atbs_core_0.spike_memory_0.n2380_o[0]\ VPWR VGND _02254_ sg13g2_buf_1
X_20859_ _02254_ _02231_ _02250_ VPWR VGND _01312_ sg13g2_mux2_1
X_20860_ \atbs_core_0.spike_memory_0.n2380_o[1]\ VPWR VGND _02255_ sg13g2_buf_1
X_20861_ _02255_ _02233_ _02250_ VPWR VGND _01313_ sg13g2_mux2_1
X_20862_ \atbs_core_0.spike_memory_0.n2360_o[3]\ VPWR VGND _02256_ sg13g2_buf_1
X_20863_ _02256_ _02073_ _02250_ VPWR VGND _01314_ sg13g2_mux2_1
X_20864_ \atbs_core_0.spike_memory_0.n2380_o[2]\ VPWR VGND _02257_ sg13g2_buf_1
X_20865_ _02257_ _02234_ _02250_ VPWR VGND _01315_ sg13g2_mux2_1
X_20866_ \atbs_core_0.spike_memory_0.n2380_o[3]\ VPWR VGND _02258_ sg13g2_buf_1
X_20867_ _02258_ _02235_ _02250_ VPWR VGND _01316_ sg13g2_mux2_1
X_20868_ \atbs_core_0.spike_memory_0.n2380_o[4]\ VPWR VGND _02259_ sg13g2_buf_1
X_20869_ _02259_ _02236_ _02250_ VPWR VGND _01317_ sg13g2_mux2_1
X_20870_ \atbs_core_0.spike_memory_0.n2380_o[5]\ VPWR VGND _02260_ sg13g2_buf_1
X_20871_ _02203_ VPWR VGND _02261_ sg13g2_buf_1
X_20872_ _02260_ _02237_ _02261_ VPWR VGND _01318_ sg13g2_mux2_1
X_20873_ \atbs_core_0.spike_memory_0.n2380_o[6]\ VPWR VGND _02262_ sg13g2_buf_1
X_20874_ _02262_ _02238_ _02261_ VPWR VGND _01319_ sg13g2_mux2_1
X_20875_ \atbs_core_0.spike_memory_0.n2380_o[7]\ VPWR VGND _02263_ sg13g2_buf_1
X_20876_ _02263_ _02240_ _02261_ VPWR VGND _01320_ sg13g2_mux2_1
X_20877_ \atbs_core_0.spike_memory_0.n2380_o[8]\ VPWR VGND _02264_ sg13g2_buf_1
X_20878_ _02264_ _02241_ _02261_ VPWR VGND _01321_ sg13g2_mux2_1
X_20879_ \atbs_core_0.spike_memory_0.n2380_o[9]\ VPWR VGND _02265_ sg13g2_buf_1
X_20880_ _02265_ _02242_ _02261_ VPWR VGND _01322_ sg13g2_mux2_1
X_20881_ \atbs_core_0.spike_memory_0.n2380_o[10]\ VPWR VGND _02266_ sg13g2_buf_1
X_20882_ _02266_ _02243_ _02261_ VPWR VGND _01323_ sg13g2_mux2_1
X_20883_ \atbs_core_0.spike_memory_0.n2380_o[11]\ VPWR VGND _02267_ sg13g2_buf_1
X_20884_ _02267_ _02245_ _02261_ VPWR VGND _01324_ sg13g2_mux2_1
X_20885_ \atbs_core_0.spike_memory_0.n2360_o[4]\ VPWR VGND _02268_ sg13g2_buf_1
X_20886_ _02268_ _02077_ _02261_ VPWR VGND _01325_ sg13g2_mux2_1
X_20887_ \atbs_core_0.spike_memory_0.n2380_o[12]\ VPWR VGND _02269_ sg13g2_buf_1
X_20888_ _02269_ _02246_ _02261_ VPWR VGND _01326_ sg13g2_mux2_1
X_20889_ \atbs_core_0.spike_memory_0.n2380_o[13]\ VPWR VGND _02270_ sg13g2_buf_1
X_20890_ _02270_ _02247_ _02261_ VPWR VGND _01327_ sg13g2_mux2_1
X_20891_ \atbs_core_0.spike_memory_0.n2380_o[14]\ VPWR VGND _02271_ sg13g2_buf_1
X_20892_ _02203_ VPWR VGND _02272_ sg13g2_buf_1
X_20893_ _02271_ _02248_ _02272_ VPWR VGND _01328_ sg13g2_mux2_1
X_20894_ \atbs_core_0.spike_memory_0.n2380_o[15]\ VPWR VGND _02273_ sg13g2_buf_1
X_20895_ _02273_ _02249_ _02272_ VPWR VGND _01329_ sg13g2_mux2_1
X_20896_ \atbs_core_0.spike_memory_0.n2380_o[16]\ VPWR VGND _02274_ sg13g2_buf_1
X_20897_ _02274_ _02251_ _02272_ VPWR VGND _01330_ sg13g2_mux2_1
X_20898_ \atbs_core_0.spike_memory_0.n2380_o[17]\ VPWR VGND _02275_ sg13g2_buf_1
X_20899_ _02275_ _02252_ _02272_ VPWR VGND _01331_ sg13g2_mux2_1
X_20900_ \atbs_core_0.spike_memory_0.n2380_o[18]\ VPWR VGND _02276_ sg13g2_buf_1
X_20901_ _02276_ _02253_ _02272_ VPWR VGND _01332_ sg13g2_mux2_1
X_20902_ \atbs_core_0.spike_memory_0.n2381_o[0]\ _02254_ _02272_ VPWR VGND _01333_ sg13g2_mux2_1
X_20903_ \atbs_core_0.spike_memory_0.n2381_o[1]\ _02255_ _02272_ VPWR VGND _01334_ sg13g2_mux2_1
X_20904_ \atbs_core_0.spike_memory_0.n2381_o[2]\ _02257_ _02272_ VPWR VGND _01335_ sg13g2_mux2_1
X_20905_ \atbs_core_0.spike_memory_0.n2360_o[5]\ VPWR VGND _02277_ sg13g2_buf_1
X_20906_ _02277_ _02082_ _02272_ VPWR VGND _01336_ sg13g2_mux2_1
X_20907_ \atbs_core_0.spike_memory_0.n2381_o[3]\ _02258_ _02272_ VPWR VGND _01337_ sg13g2_mux2_1
X_20908_ _02074_ VPWR VGND _02278_ sg13g2_buf_1
X_20909_ _02278_ VPWR VGND _02279_ sg13g2_buf_1
X_20910_ \atbs_core_0.spike_memory_0.n2381_o[4]\ _02259_ _02279_ VPWR VGND _01338_ sg13g2_mux2_1
X_20911_ \atbs_core_0.spike_memory_0.n2381_o[5]\ _02260_ _02279_ VPWR VGND _01339_ sg13g2_mux2_1
X_20912_ \atbs_core_0.spike_memory_0.n2381_o[6]\ _02262_ _02279_ VPWR VGND _01340_ sg13g2_mux2_1
X_20913_ \atbs_core_0.spike_memory_0.n2381_o[7]\ _02263_ _02279_ VPWR VGND _01341_ sg13g2_mux2_1
X_20914_ \atbs_core_0.spike_memory_0.n2381_o[8]\ _02264_ _02279_ VPWR VGND _01342_ sg13g2_mux2_1
X_20915_ \atbs_core_0.spike_memory_0.n2381_o[9]\ _02265_ _02279_ VPWR VGND _01343_ sg13g2_mux2_1
X_20916_ \atbs_core_0.spike_memory_0.n2381_o[10]\ _02266_ _02279_ VPWR VGND _01344_ sg13g2_mux2_1
X_20917_ \atbs_core_0.spike_memory_0.n2381_o[11]\ _02267_ _02279_ VPWR VGND _01345_ sg13g2_mux2_1
X_20918_ \atbs_core_0.spike_memory_0.n2381_o[12]\ _02269_ _02279_ VPWR VGND _01346_ sg13g2_mux2_1
X_20919_ \atbs_core_0.spike_memory_0.n2360_o[6]\ VPWR VGND _02280_ sg13g2_buf_1
X_20920_ _02280_ _02094_ _02279_ VPWR VGND _01347_ sg13g2_mux2_1
X_20921_ _02278_ VPWR VGND _02281_ sg13g2_buf_1
X_20922_ \atbs_core_0.spike_memory_0.n2381_o[13]\ _02270_ _02281_ VPWR VGND _01348_ sg13g2_mux2_1
X_20923_ \atbs_core_0.spike_memory_0.n2381_o[14]\ _02271_ _02281_ VPWR VGND _01349_ sg13g2_mux2_1
X_20924_ \atbs_core_0.spike_memory_0.n2381_o[15]\ _02273_ _02281_ VPWR VGND _01350_ sg13g2_mux2_1
X_20925_ \atbs_core_0.spike_memory_0.n2381_o[16]\ _02274_ _02281_ VPWR VGND _01351_ sg13g2_mux2_1
X_20926_ \atbs_core_0.spike_memory_0.n2381_o[17]\ _02275_ _02281_ VPWR VGND _01352_ sg13g2_mux2_1
X_20927_ \atbs_core_0.spike_memory_0.n2381_o[18]\ _02276_ _02281_ VPWR VGND _01353_ sg13g2_mux2_1
X_20928_ \atbs_core_0.spike_memory_0.n2382_o[0]\ \atbs_core_0.spike_memory_0.n2381_o[0]\ _02281_ VPWR VGND _01354_ sg13g2_mux2_1
X_20929_ \atbs_core_0.spike_memory_0.n2382_o[1]\ \atbs_core_0.spike_memory_0.n2381_o[1]\ _02281_ VPWR VGND _01355_ sg13g2_mux2_1
X_20930_ \atbs_core_0.spike_memory_0.n2382_o[2]\ \atbs_core_0.spike_memory_0.n2381_o[2]\ _02281_ VPWR VGND _01356_ sg13g2_mux2_1
X_20931_ \atbs_core_0.spike_memory_0.n2382_o[3]\ \atbs_core_0.spike_memory_0.n2381_o[3]\ _02281_ VPWR VGND _01357_ sg13g2_mux2_1
X_20932_ \atbs_core_0.spike_memory_0.n2360_o[7]\ VPWR VGND _02282_ sg13g2_buf_1
X_20933_ _02278_ VPWR VGND _02283_ sg13g2_buf_1
X_20934_ _02282_ _02106_ _02283_ VPWR VGND _01358_ sg13g2_mux2_1
X_20935_ \atbs_core_0.spike_memory_0.n2382_o[4]\ \atbs_core_0.spike_memory_0.n2381_o[4]\ _02283_ VPWR VGND _01359_ sg13g2_mux2_1
X_20936_ \atbs_core_0.spike_memory_0.n2382_o[5]\ \atbs_core_0.spike_memory_0.n2381_o[5]\ _02283_ VPWR VGND _01360_ sg13g2_mux2_1
X_20937_ \atbs_core_0.spike_memory_0.n2382_o[6]\ \atbs_core_0.spike_memory_0.n2381_o[6]\ _02283_ VPWR VGND _01361_ sg13g2_mux2_1
X_20938_ \atbs_core_0.spike_memory_0.n2382_o[7]\ \atbs_core_0.spike_memory_0.n2381_o[7]\ _02283_ VPWR VGND _01362_ sg13g2_mux2_1
X_20939_ \atbs_core_0.spike_memory_0.n2382_o[8]\ \atbs_core_0.spike_memory_0.n2381_o[8]\ _02283_ VPWR VGND _01363_ sg13g2_mux2_1
X_20940_ \atbs_core_0.spike_memory_0.n2382_o[9]\ \atbs_core_0.spike_memory_0.n2381_o[9]\ _02283_ VPWR VGND _01364_ sg13g2_mux2_1
X_20941_ \atbs_core_0.spike_memory_0.n2382_o[10]\ \atbs_core_0.spike_memory_0.n2381_o[10]\ _02283_ VPWR VGND _01365_ sg13g2_mux2_1
X_20942_ \atbs_core_0.spike_memory_0.n2382_o[11]\ \atbs_core_0.spike_memory_0.n2381_o[11]\ _02283_ VPWR VGND _01366_ sg13g2_mux2_1
X_20943_ \atbs_core_0.spike_memory_0.n2382_o[12]\ \atbs_core_0.spike_memory_0.n2381_o[12]\ _02283_ VPWR VGND _01367_ sg13g2_mux2_1
X_20944_ _02278_ VPWR VGND _02284_ sg13g2_buf_1
X_20945_ \atbs_core_0.spike_memory_0.n2382_o[13]\ \atbs_core_0.spike_memory_0.n2381_o[13]\ _02284_ VPWR VGND _01368_ sg13g2_mux2_1
X_20946_ \atbs_core_0.spike_memory_0.n2360_o[8]\ VPWR VGND _02285_ sg13g2_buf_1
X_20947_ _02285_ _02118_ _02284_ VPWR VGND _01369_ sg13g2_mux2_1
X_20948_ \atbs_core_0.spike_memory_0.n2382_o[14]\ \atbs_core_0.spike_memory_0.n2381_o[14]\ _02284_ VPWR VGND _01370_ sg13g2_mux2_1
X_20949_ \atbs_core_0.spike_memory_0.n2382_o[15]\ \atbs_core_0.spike_memory_0.n2381_o[15]\ _02284_ VPWR VGND _01371_ sg13g2_mux2_1
X_20950_ \atbs_core_0.spike_memory_0.n2382_o[16]\ \atbs_core_0.spike_memory_0.n2381_o[16]\ _02284_ VPWR VGND _01372_ sg13g2_mux2_1
X_20951_ \atbs_core_0.spike_memory_0.n2382_o[17]\ \atbs_core_0.spike_memory_0.n2381_o[17]\ _02284_ VPWR VGND _01373_ sg13g2_mux2_1
X_20952_ \atbs_core_0.spike_memory_0.n2382_o[18]\ \atbs_core_0.spike_memory_0.n2381_o[18]\ _02284_ VPWR VGND _01374_ sg13g2_mux2_1
X_20953_ \atbs_core_0.spike_memory_0.n2383_o[0]\ VPWR VGND _02286_ sg13g2_buf_1
X_20954_ _02286_ \atbs_core_0.spike_memory_0.n2382_o[0]\ _02284_ VPWR VGND _01375_ sg13g2_mux2_1
X_20955_ \atbs_core_0.spike_memory_0.n2383_o[1]\ VPWR VGND _02287_ sg13g2_buf_1
X_20956_ _02287_ \atbs_core_0.spike_memory_0.n2382_o[1]\ _02284_ VPWR VGND _01376_ sg13g2_mux2_1
X_20957_ \atbs_core_0.spike_memory_0.n2383_o[2]\ VPWR VGND _02288_ sg13g2_buf_1
X_20958_ _02288_ \atbs_core_0.spike_memory_0.n2382_o[2]\ _02284_ VPWR VGND _01377_ sg13g2_mux2_1
X_20959_ \atbs_core_0.spike_memory_0.n2383_o[3]\ VPWR VGND _02289_ sg13g2_buf_1
X_20960_ _02278_ VPWR VGND _02290_ sg13g2_buf_1
X_20961_ _02289_ \atbs_core_0.spike_memory_0.n2382_o[3]\ _02290_ VPWR VGND _01378_ sg13g2_mux2_1
X_20962_ \atbs_core_0.spike_memory_0.n2383_o[4]\ VPWR VGND _02291_ sg13g2_buf_1
X_20963_ _02291_ \atbs_core_0.spike_memory_0.n2382_o[4]\ _02290_ VPWR VGND _01379_ sg13g2_mux2_1
X_20964_ \atbs_core_0.spike_memory_0.n2360_o[9]\ VPWR VGND _02292_ sg13g2_buf_1
X_20965_ _02292_ _02125_ _02290_ VPWR VGND _01380_ sg13g2_mux2_1
X_20966_ \atbs_core_0.spike_memory_0.n2383_o[5]\ VPWR VGND _02293_ sg13g2_buf_1
X_20967_ _02293_ \atbs_core_0.spike_memory_0.n2382_o[5]\ _02290_ VPWR VGND _01381_ sg13g2_mux2_1
X_20968_ \atbs_core_0.spike_memory_0.n2383_o[6]\ VPWR VGND _02294_ sg13g2_buf_1
X_20969_ _02294_ \atbs_core_0.spike_memory_0.n2382_o[6]\ _02290_ VPWR VGND _01382_ sg13g2_mux2_1
X_20970_ \atbs_core_0.spike_memory_0.n2383_o[7]\ VPWR VGND _02295_ sg13g2_buf_1
X_20971_ _02295_ \atbs_core_0.spike_memory_0.n2382_o[7]\ _02290_ VPWR VGND _01383_ sg13g2_mux2_1
X_20972_ \atbs_core_0.spike_memory_0.n2383_o[8]\ VPWR VGND _02296_ sg13g2_buf_1
X_20973_ _02296_ \atbs_core_0.spike_memory_0.n2382_o[8]\ _02290_ VPWR VGND _01384_ sg13g2_mux2_1
X_20974_ \atbs_core_0.spike_memory_0.n2383_o[9]\ VPWR VGND _02297_ sg13g2_buf_1
X_20975_ _02297_ \atbs_core_0.spike_memory_0.n2382_o[9]\ _02290_ VPWR VGND _01385_ sg13g2_mux2_1
X_20976_ \atbs_core_0.spike_memory_0.n2383_o[10]\ VPWR VGND _02298_ sg13g2_buf_1
X_20977_ _02298_ \atbs_core_0.spike_memory_0.n2382_o[10]\ _02290_ VPWR VGND _01386_ sg13g2_mux2_1
X_20978_ \atbs_core_0.spike_memory_0.n2383_o[11]\ VPWR VGND _02299_ sg13g2_buf_1
X_20979_ _02299_ \atbs_core_0.spike_memory_0.n2382_o[11]\ _02290_ VPWR VGND _01387_ sg13g2_mux2_1
X_20980_ \atbs_core_0.spike_memory_0.n2383_o[12]\ VPWR VGND _02300_ sg13g2_buf_1
X_20981_ _02278_ VPWR VGND _02301_ sg13g2_buf_1
X_20982_ _02300_ \atbs_core_0.spike_memory_0.n2382_o[12]\ _02301_ VPWR VGND _01388_ sg13g2_mux2_1
X_20983_ \atbs_core_0.spike_memory_0.n2383_o[13]\ VPWR VGND _02302_ sg13g2_buf_1
X_20984_ _02302_ \atbs_core_0.spike_memory_0.n2382_o[13]\ _02301_ VPWR VGND _01389_ sg13g2_mux2_1
X_20985_ \atbs_core_0.spike_memory_0.n2383_o[14]\ VPWR VGND _02303_ sg13g2_buf_1
X_20986_ _02303_ \atbs_core_0.spike_memory_0.n2382_o[14]\ _02301_ VPWR VGND _01390_ sg13g2_mux2_1
X_20987_ \atbs_core_0.spike_memory_0.n2360_o[10]\ VPWR VGND _02304_ sg13g2_buf_1
X_20988_ _02304_ _02129_ _02301_ VPWR VGND _01391_ sg13g2_mux2_1
X_20989_ \atbs_core_0.spike_memory_0.n2383_o[15]\ VPWR VGND _02305_ sg13g2_buf_1
X_20990_ _02305_ \atbs_core_0.spike_memory_0.n2382_o[15]\ _02301_ VPWR VGND _01392_ sg13g2_mux2_1
X_20991_ \atbs_core_0.spike_memory_0.n2383_o[16]\ VPWR VGND _02306_ sg13g2_buf_1
X_20992_ _02306_ \atbs_core_0.spike_memory_0.n2382_o[16]\ _02301_ VPWR VGND _01393_ sg13g2_mux2_1
X_20993_ \atbs_core_0.spike_memory_0.n2383_o[17]\ VPWR VGND _02307_ sg13g2_buf_1
X_20994_ _02307_ \atbs_core_0.spike_memory_0.n2382_o[17]\ _02301_ VPWR VGND _01394_ sg13g2_mux2_1
X_20995_ \atbs_core_0.spike_memory_0.n2383_o[18]\ VPWR VGND _02308_ sg13g2_buf_1
X_20996_ _02308_ \atbs_core_0.spike_memory_0.n2382_o[18]\ _02301_ VPWR VGND _01395_ sg13g2_mux2_1
X_20997_ \atbs_core_0.spike_memory_0.n2384_o[0]\ VPWR VGND _02309_ sg13g2_buf_1
X_20998_ _02309_ _02286_ _02301_ VPWR VGND _01396_ sg13g2_mux2_1
X_20999_ \atbs_core_0.spike_memory_0.n2384_o[1]\ VPWR VGND _02310_ sg13g2_buf_1
X_21000_ _02310_ _02287_ _02301_ VPWR VGND _01397_ sg13g2_mux2_1
X_21001_ \atbs_core_0.spike_memory_0.n2384_o[2]\ VPWR VGND _02311_ sg13g2_buf_1
X_21002_ _02278_ VPWR VGND _02312_ sg13g2_buf_1
X_21003_ _02311_ _02288_ _02312_ VPWR VGND _01398_ sg13g2_mux2_1
X_21004_ \atbs_core_0.spike_memory_0.n2384_o[3]\ VPWR VGND _02313_ sg13g2_buf_1
X_21005_ _02313_ _02289_ _02312_ VPWR VGND _01399_ sg13g2_mux2_1
X_21006_ \atbs_core_0.spike_memory_0.n2384_o[4]\ VPWR VGND _02314_ sg13g2_buf_1
X_21007_ _02314_ _02291_ _02312_ VPWR VGND _01400_ sg13g2_mux2_1
X_21008_ \atbs_core_0.spike_memory_0.n2384_o[5]\ VPWR VGND _02315_ sg13g2_buf_1
X_21009_ _02315_ _02293_ _02312_ VPWR VGND _01401_ sg13g2_mux2_1
X_21010_ \atbs_core_0.spike_memory_0.n2360_o[11]\ VPWR VGND _02316_ sg13g2_buf_1
X_21011_ _02316_ _02131_ _02312_ VPWR VGND _01402_ sg13g2_mux2_1
X_21012_ \atbs_core_0.spike_memory_0.n2358_o[4]\ \atbs_core_0.spike_memory_0.a_data[4]\ _02312_ VPWR VGND _01403_ sg13g2_mux2_1
X_21013_ \atbs_core_0.spike_memory_0.n2384_o[6]\ VPWR VGND _02317_ sg13g2_buf_1
X_21014_ _02317_ _02294_ _02312_ VPWR VGND _01404_ sg13g2_mux2_1
X_21015_ \atbs_core_0.spike_memory_0.n2384_o[7]\ VPWR VGND _02318_ sg13g2_buf_1
X_21016_ _02318_ _02295_ _02312_ VPWR VGND _01405_ sg13g2_mux2_1
X_21017_ \atbs_core_0.spike_memory_0.n2384_o[8]\ VPWR VGND _02319_ sg13g2_buf_1
X_21018_ _02319_ _02296_ _02312_ VPWR VGND _01406_ sg13g2_mux2_1
X_21019_ \atbs_core_0.spike_memory_0.n2384_o[9]\ VPWR VGND _02320_ sg13g2_buf_1
X_21020_ _02320_ _02297_ _02312_ VPWR VGND _01407_ sg13g2_mux2_1
X_21021_ \atbs_core_0.spike_memory_0.n2384_o[10]\ VPWR VGND _02321_ sg13g2_buf_1
X_21022_ _02074_ VPWR VGND _02322_ sg13g2_buf_1
X_21023_ _02322_ VPWR VGND _02323_ sg13g2_buf_1
X_21024_ _02321_ _02298_ _02323_ VPWR VGND _01408_ sg13g2_mux2_1
X_21025_ \atbs_core_0.spike_memory_0.n2384_o[11]\ VPWR VGND _02324_ sg13g2_buf_1
X_21026_ _02324_ _02299_ _02323_ VPWR VGND _01409_ sg13g2_mux2_1
X_21027_ \atbs_core_0.spike_memory_0.n2384_o[12]\ VPWR VGND _02325_ sg13g2_buf_1
X_21028_ _02325_ _02300_ _02323_ VPWR VGND _01410_ sg13g2_mux2_1
X_21029_ \atbs_core_0.spike_memory_0.n2384_o[13]\ VPWR VGND _02326_ sg13g2_buf_1
X_21030_ _02326_ _02302_ _02323_ VPWR VGND _01411_ sg13g2_mux2_1
X_21031_ \atbs_core_0.spike_memory_0.n2384_o[14]\ VPWR VGND _02327_ sg13g2_buf_1
X_21032_ _02327_ _02303_ _02323_ VPWR VGND _01412_ sg13g2_mux2_1
X_21033_ \atbs_core_0.spike_memory_0.n2384_o[15]\ VPWR VGND _02328_ sg13g2_buf_1
X_21034_ _02328_ _02305_ _02323_ VPWR VGND _01413_ sg13g2_mux2_1
X_21035_ \atbs_core_0.spike_memory_0.n2360_o[12]\ VPWR VGND _02329_ sg13g2_buf_1
X_21036_ _02329_ _02133_ _02323_ VPWR VGND _01414_ sg13g2_mux2_1
X_21037_ \atbs_core_0.spike_memory_0.n2384_o[16]\ VPWR VGND _02330_ sg13g2_buf_1
X_21038_ _02330_ _02306_ _02323_ VPWR VGND _01415_ sg13g2_mux2_1
X_21039_ \atbs_core_0.spike_memory_0.n2384_o[17]\ VPWR VGND _02331_ sg13g2_buf_1
X_21040_ _02331_ _02307_ _02323_ VPWR VGND _01416_ sg13g2_mux2_1
X_21041_ \atbs_core_0.spike_memory_0.n2384_o[18]\ VPWR VGND _02332_ sg13g2_buf_1
X_21042_ _02332_ _02308_ _02323_ VPWR VGND _01417_ sg13g2_mux2_1
X_21043_ _02322_ VPWR VGND _02333_ sg13g2_buf_1
X_21044_ \atbs_core_0.spike_memory_0.n2385_o[0]\ _02309_ _02333_ VPWR VGND _01418_ sg13g2_mux2_1
X_21045_ \atbs_core_0.spike_memory_0.n2385_o[1]\ _02310_ _02333_ VPWR VGND _01419_ sg13g2_mux2_1
X_21046_ \atbs_core_0.spike_memory_0.n2385_o[2]\ _02311_ _02333_ VPWR VGND _01420_ sg13g2_mux2_1
X_21047_ \atbs_core_0.spike_memory_0.n2385_o[3]\ _02313_ _02333_ VPWR VGND _01421_ sg13g2_mux2_1
X_21048_ \atbs_core_0.spike_memory_0.n2385_o[4]\ _02314_ _02333_ VPWR VGND _01422_ sg13g2_mux2_1
X_21049_ \atbs_core_0.spike_memory_0.n2385_o[5]\ _02315_ _02333_ VPWR VGND _01423_ sg13g2_mux2_1
X_21050_ \atbs_core_0.spike_memory_0.n2385_o[6]\ _02317_ _02333_ VPWR VGND _01424_ sg13g2_mux2_1
X_21051_ \atbs_core_0.spike_memory_0.n2360_o[13]\ VPWR VGND _02334_ sg13g2_buf_1
X_21052_ _02334_ _02142_ _02333_ VPWR VGND _01425_ sg13g2_mux2_1
X_21053_ \atbs_core_0.spike_memory_0.n2385_o[7]\ _02318_ _02333_ VPWR VGND _01426_ sg13g2_mux2_1
X_21054_ \atbs_core_0.spike_memory_0.n2385_o[8]\ _02319_ _02333_ VPWR VGND _01427_ sg13g2_mux2_1
X_21055_ _02322_ VPWR VGND _02335_ sg13g2_buf_1
X_21056_ \atbs_core_0.spike_memory_0.n2385_o[9]\ _02320_ _02335_ VPWR VGND _01428_ sg13g2_mux2_1
X_21057_ \atbs_core_0.spike_memory_0.n2385_o[10]\ _02321_ _02335_ VPWR VGND _01429_ sg13g2_mux2_1
X_21058_ \atbs_core_0.spike_memory_0.n2385_o[11]\ _02324_ _02335_ VPWR VGND _01430_ sg13g2_mux2_1
X_21059_ \atbs_core_0.spike_memory_0.n2385_o[12]\ _02325_ _02335_ VPWR VGND _01431_ sg13g2_mux2_1
X_21060_ \atbs_core_0.spike_memory_0.n2385_o[13]\ _02326_ _02335_ VPWR VGND _01432_ sg13g2_mux2_1
X_21061_ \atbs_core_0.spike_memory_0.n2385_o[14]\ _02327_ _02335_ VPWR VGND _01433_ sg13g2_mux2_1
X_21062_ \atbs_core_0.spike_memory_0.n2385_o[15]\ _02328_ _02335_ VPWR VGND _01434_ sg13g2_mux2_1
X_21063_ \atbs_core_0.spike_memory_0.n2385_o[16]\ _02330_ _02335_ VPWR VGND _01435_ sg13g2_mux2_1
X_21064_ \atbs_core_0.spike_memory_0.n2360_o[14]\ VPWR VGND _02336_ sg13g2_buf_1
X_21065_ _02336_ _02154_ _02335_ VPWR VGND _01436_ sg13g2_mux2_1
X_21066_ \atbs_core_0.spike_memory_0.n2385_o[17]\ _02331_ _02335_ VPWR VGND _01437_ sg13g2_mux2_1
X_21067_ _02322_ VPWR VGND _02337_ sg13g2_buf_1
X_21068_ \atbs_core_0.spike_memory_0.n2385_o[18]\ _02332_ _02337_ VPWR VGND _01438_ sg13g2_mux2_1
X_21069_ \atbs_core_0.spike_memory_0.n2386_o[0]\ \atbs_core_0.spike_memory_0.n2385_o[0]\ _02337_ VPWR VGND _01439_ sg13g2_mux2_1
X_21070_ \atbs_core_0.spike_memory_0.n2386_o[1]\ \atbs_core_0.spike_memory_0.n2385_o[1]\ _02337_ VPWR VGND _01440_ sg13g2_mux2_1
X_21071_ \atbs_core_0.spike_memory_0.n2386_o[2]\ \atbs_core_0.spike_memory_0.n2385_o[2]\ _02337_ VPWR VGND _01441_ sg13g2_mux2_1
X_21072_ \atbs_core_0.spike_memory_0.n2386_o[3]\ \atbs_core_0.spike_memory_0.n2385_o[3]\ _02337_ VPWR VGND _01442_ sg13g2_mux2_1
X_21073_ \atbs_core_0.spike_memory_0.n2386_o[4]\ \atbs_core_0.spike_memory_0.n2385_o[4]\ _02337_ VPWR VGND _01443_ sg13g2_mux2_1
X_21074_ \atbs_core_0.spike_memory_0.n2386_o[5]\ \atbs_core_0.spike_memory_0.n2385_o[5]\ _02337_ VPWR VGND _01444_ sg13g2_mux2_1
X_21075_ \atbs_core_0.spike_memory_0.n2386_o[6]\ \atbs_core_0.spike_memory_0.n2385_o[6]\ _02337_ VPWR VGND _01445_ sg13g2_mux2_1
X_21076_ \atbs_core_0.spike_memory_0.n2386_o[7]\ \atbs_core_0.spike_memory_0.n2385_o[7]\ _02337_ VPWR VGND _01446_ sg13g2_mux2_1
X_21077_ \atbs_core_0.spike_memory_0.n2360_o[15]\ VPWR VGND _02338_ sg13g2_buf_1
X_21078_ _02338_ _02166_ _02337_ VPWR VGND _01447_ sg13g2_mux2_1
X_21079_ _02322_ VPWR VGND _02339_ sg13g2_buf_1
X_21080_ \atbs_core_0.spike_memory_0.n2386_o[8]\ \atbs_core_0.spike_memory_0.n2385_o[8]\ _02339_ VPWR VGND _01448_ sg13g2_mux2_1
X_21081_ \atbs_core_0.spike_memory_0.n2386_o[9]\ \atbs_core_0.spike_memory_0.n2385_o[9]\ _02339_ VPWR VGND _01449_ sg13g2_mux2_1
X_21082_ \atbs_core_0.spike_memory_0.n2386_o[10]\ \atbs_core_0.spike_memory_0.n2385_o[10]\ _02339_ VPWR VGND _01450_ sg13g2_mux2_1
X_21083_ \atbs_core_0.spike_memory_0.n2386_o[11]\ \atbs_core_0.spike_memory_0.n2385_o[11]\ _02339_ VPWR VGND _01451_ sg13g2_mux2_1
X_21084_ \atbs_core_0.spike_memory_0.n2386_o[12]\ \atbs_core_0.spike_memory_0.n2385_o[12]\ _02339_ VPWR VGND _01452_ sg13g2_mux2_1
X_21085_ \atbs_core_0.spike_memory_0.n2386_o[13]\ \atbs_core_0.spike_memory_0.n2385_o[13]\ _02339_ VPWR VGND _01453_ sg13g2_mux2_1
X_21086_ \atbs_core_0.spike_memory_0.n2386_o[14]\ \atbs_core_0.spike_memory_0.n2385_o[14]\ _02339_ VPWR VGND _01454_ sg13g2_mux2_1
X_21087_ \atbs_core_0.spike_memory_0.n2386_o[15]\ \atbs_core_0.spike_memory_0.n2385_o[15]\ _02339_ VPWR VGND _01455_ sg13g2_mux2_1
X_21088_ \atbs_core_0.spike_memory_0.n2386_o[16]\ \atbs_core_0.spike_memory_0.n2385_o[16]\ _02339_ VPWR VGND _01456_ sg13g2_mux2_1
X_21089_ \atbs_core_0.spike_memory_0.n2386_o[17]\ \atbs_core_0.spike_memory_0.n2385_o[17]\ _02339_ VPWR VGND _01457_ sg13g2_mux2_1
X_21090_ \atbs_core_0.spike_memory_0.n2360_o[16]\ VPWR VGND _02340_ sg13g2_buf_1
X_21091_ _02322_ VPWR VGND _02341_ sg13g2_buf_1
X_21092_ _02340_ _02178_ _02341_ VPWR VGND _01458_ sg13g2_mux2_1
X_21093_ \atbs_core_0.spike_memory_0.n2386_o[18]\ \atbs_core_0.spike_memory_0.n2385_o[18]\ _02341_ VPWR VGND _01459_ sg13g2_mux2_1
X_21094_ \atbs_core_0.spike_memory_0.n2387_o[0]\ VPWR VGND _02342_ sg13g2_buf_1
X_21095_ _02342_ \atbs_core_0.spike_memory_0.n2386_o[0]\ _02341_ VPWR VGND _01460_ sg13g2_mux2_1
X_21096_ \atbs_core_0.spike_memory_0.n2387_o[1]\ VPWR VGND _02343_ sg13g2_buf_1
X_21097_ _02343_ \atbs_core_0.spike_memory_0.n2386_o[1]\ _02341_ VPWR VGND _01461_ sg13g2_mux2_1
X_21098_ \atbs_core_0.spike_memory_0.n2387_o[2]\ VPWR VGND _02344_ sg13g2_buf_1
X_21099_ _02344_ \atbs_core_0.spike_memory_0.n2386_o[2]\ _02341_ VPWR VGND _01462_ sg13g2_mux2_1
X_21100_ \atbs_core_0.spike_memory_0.n2387_o[3]\ VPWR VGND _02345_ sg13g2_buf_1
X_21101_ _02345_ \atbs_core_0.spike_memory_0.n2386_o[3]\ _02341_ VPWR VGND _01463_ sg13g2_mux2_1
X_21102_ \atbs_core_0.spike_memory_0.n2387_o[4]\ VPWR VGND _02346_ sg13g2_buf_1
X_21103_ _02346_ \atbs_core_0.spike_memory_0.n2386_o[4]\ _02341_ VPWR VGND _01464_ sg13g2_mux2_1
X_21104_ \atbs_core_0.spike_memory_0.n2387_o[5]\ VPWR VGND _02347_ sg13g2_buf_1
X_21105_ _02347_ \atbs_core_0.spike_memory_0.n2386_o[5]\ _02341_ VPWR VGND _01465_ sg13g2_mux2_1
X_21106_ \atbs_core_0.spike_memory_0.n2387_o[6]\ VPWR VGND _02348_ sg13g2_buf_1
X_21107_ _02348_ \atbs_core_0.spike_memory_0.n2386_o[6]\ _02341_ VPWR VGND _01466_ sg13g2_mux2_1
X_21108_ \atbs_core_0.spike_memory_0.n2387_o[7]\ VPWR VGND _02349_ sg13g2_buf_1
X_21109_ _02349_ \atbs_core_0.spike_memory_0.n2386_o[7]\ _02341_ VPWR VGND _01467_ sg13g2_mux2_1
X_21110_ \atbs_core_0.spike_memory_0.n2387_o[8]\ VPWR VGND _02350_ sg13g2_buf_1
X_21111_ _02322_ VPWR VGND _02351_ sg13g2_buf_1
X_21112_ _02350_ \atbs_core_0.spike_memory_0.n2386_o[8]\ _02351_ VPWR VGND _01468_ sg13g2_mux2_1
X_21113_ \atbs_core_0.spike_memory_0.n2360_o[17]\ VPWR VGND _02352_ sg13g2_buf_1
X_21114_ _02352_ _02202_ _02351_ VPWR VGND _01469_ sg13g2_mux2_1
X_21115_ \atbs_core_0.spike_memory_0.n2387_o[9]\ VPWR VGND _02353_ sg13g2_buf_1
X_21116_ _02353_ \atbs_core_0.spike_memory_0.n2386_o[9]\ _02351_ VPWR VGND _01470_ sg13g2_mux2_1
X_21117_ \atbs_core_0.spike_memory_0.n2387_o[10]\ VPWR VGND _02354_ sg13g2_buf_1
X_21118_ _02354_ \atbs_core_0.spike_memory_0.n2386_o[10]\ _02351_ VPWR VGND _01471_ sg13g2_mux2_1
X_21119_ \atbs_core_0.spike_memory_0.n2387_o[11]\ VPWR VGND _02355_ sg13g2_buf_1
X_21120_ _02355_ \atbs_core_0.spike_memory_0.n2386_o[11]\ _02351_ VPWR VGND _01472_ sg13g2_mux2_1
X_21121_ \atbs_core_0.spike_memory_0.n2387_o[12]\ VPWR VGND _02356_ sg13g2_buf_1
X_21122_ _02356_ \atbs_core_0.spike_memory_0.n2386_o[12]\ _02351_ VPWR VGND _01473_ sg13g2_mux2_1
X_21123_ \atbs_core_0.spike_memory_0.n2387_o[13]\ VPWR VGND _02357_ sg13g2_buf_1
X_21124_ _02357_ \atbs_core_0.spike_memory_0.n2386_o[13]\ _02351_ VPWR VGND _01474_ sg13g2_mux2_1
X_21125_ \atbs_core_0.spike_memory_0.n2387_o[14]\ VPWR VGND _02358_ sg13g2_buf_1
X_21126_ _02358_ \atbs_core_0.spike_memory_0.n2386_o[14]\ _02351_ VPWR VGND _01475_ sg13g2_mux2_1
X_21127_ \atbs_core_0.spike_memory_0.n2387_o[15]\ VPWR VGND _02359_ sg13g2_buf_1
X_21128_ _02359_ \atbs_core_0.spike_memory_0.n2386_o[15]\ _02351_ VPWR VGND _01476_ sg13g2_mux2_1
X_21129_ \atbs_core_0.spike_memory_0.n2387_o[16]\ VPWR VGND _02360_ sg13g2_buf_1
X_21130_ _02360_ \atbs_core_0.spike_memory_0.n2386_o[16]\ _02351_ VPWR VGND _01477_ sg13g2_mux2_1
X_21131_ \atbs_core_0.spike_memory_0.n2387_o[17]\ VPWR VGND _02361_ sg13g2_buf_1
X_21132_ _02074_ VPWR VGND _02362_ sg13g2_buf_1
X_21133_ _02362_ VPWR VGND _02363_ sg13g2_buf_1
X_21134_ _02361_ \atbs_core_0.spike_memory_0.n2386_o[17]\ _02363_ VPWR VGND _01478_ sg13g2_mux2_1
X_21135_ \atbs_core_0.spike_memory_0.n2387_o[18]\ VPWR VGND _02364_ sg13g2_buf_1
X_21136_ _02364_ \atbs_core_0.spike_memory_0.n2386_o[18]\ _02363_ VPWR VGND _01479_ sg13g2_mux2_1
X_21137_ \atbs_core_0.spike_memory_0.n2360_o[18]\ VPWR VGND _02365_ sg13g2_buf_1
X_21138_ _02365_ _02227_ _02363_ VPWR VGND _01480_ sg13g2_mux2_1
X_21139_ \atbs_core_0.spike_memory_0.n2388_o[0]\ VPWR VGND _02366_ sg13g2_buf_1
X_21140_ _02366_ _02342_ _02363_ VPWR VGND _01481_ sg13g2_mux2_1
X_21141_ \atbs_core_0.spike_memory_0.n2388_o[1]\ VPWR VGND _02367_ sg13g2_buf_1
X_21142_ _02367_ _02343_ _02363_ VPWR VGND _01482_ sg13g2_mux2_1
X_21143_ \atbs_core_0.spike_memory_0.n2388_o[2]\ VPWR VGND _02368_ sg13g2_buf_1
X_21144_ _02368_ _02344_ _02363_ VPWR VGND _01483_ sg13g2_mux2_1
X_21145_ \atbs_core_0.spike_memory_0.n2388_o[3]\ VPWR VGND _02369_ sg13g2_buf_1
X_21146_ _02369_ _02345_ _02363_ VPWR VGND _01484_ sg13g2_mux2_1
X_21147_ \atbs_core_0.spike_memory_0.n2388_o[4]\ VPWR VGND _02370_ sg13g2_buf_1
X_21148_ _02370_ _02346_ _02363_ VPWR VGND _01485_ sg13g2_mux2_1
X_21149_ \atbs_core_0.spike_memory_0.n2388_o[5]\ VPWR VGND _02371_ sg13g2_buf_1
X_21150_ _02371_ _02347_ _02363_ VPWR VGND _01486_ sg13g2_mux2_1
X_21151_ \atbs_core_0.spike_memory_0.n2388_o[6]\ VPWR VGND _02372_ sg13g2_buf_1
X_21152_ _02372_ _02348_ _02363_ VPWR VGND _01487_ sg13g2_mux2_1
X_21153_ \atbs_core_0.spike_memory_0.n2388_o[7]\ VPWR VGND _02373_ sg13g2_buf_1
X_21154_ _02362_ VPWR VGND _02374_ sg13g2_buf_1
X_21155_ _02373_ _02349_ _02374_ VPWR VGND _01488_ sg13g2_mux2_1
X_21156_ \atbs_core_0.spike_memory_0.n2388_o[8]\ VPWR VGND _02375_ sg13g2_buf_1
X_21157_ _02375_ _02350_ _02374_ VPWR VGND _01489_ sg13g2_mux2_1
X_21158_ \atbs_core_0.spike_memory_0.n2388_o[9]\ VPWR VGND _02376_ sg13g2_buf_1
X_21159_ _02376_ _02353_ _02374_ VPWR VGND _01490_ sg13g2_mux2_1
X_21160_ \atbs_core_0.spike_memory_0.n2361_o[0]\ _02229_ _02374_ VPWR VGND _01491_ sg13g2_mux2_1
X_21161_ \atbs_core_0.spike_memory_0.n2388_o[10]\ VPWR VGND _02377_ sg13g2_buf_1
X_21162_ _02377_ _02354_ _02374_ VPWR VGND _01492_ sg13g2_mux2_1
X_21163_ \atbs_core_0.spike_memory_0.n2388_o[11]\ VPWR VGND _02378_ sg13g2_buf_1
X_21164_ _02378_ _02355_ _02374_ VPWR VGND _01493_ sg13g2_mux2_1
X_21165_ \atbs_core_0.spike_memory_0.n2388_o[12]\ VPWR VGND _02379_ sg13g2_buf_1
X_21166_ _02379_ _02356_ _02374_ VPWR VGND _01494_ sg13g2_mux2_1
X_21167_ \atbs_core_0.spike_memory_0.n2388_o[13]\ VPWR VGND _02380_ sg13g2_buf_1
X_21168_ _02380_ _02357_ _02374_ VPWR VGND _01495_ sg13g2_mux2_1
X_21169_ \atbs_core_0.spike_memory_0.n2388_o[14]\ VPWR VGND _02381_ sg13g2_buf_1
X_21170_ _02381_ _02358_ _02374_ VPWR VGND _01496_ sg13g2_mux2_1
X_21171_ \atbs_core_0.spike_memory_0.n2388_o[15]\ VPWR VGND _02382_ sg13g2_buf_1
X_21172_ _02382_ _02359_ _02374_ VPWR VGND _01497_ sg13g2_mux2_1
X_21173_ \atbs_core_0.spike_memory_0.n2388_o[16]\ VPWR VGND _02383_ sg13g2_buf_1
X_21174_ _02362_ VPWR VGND _02384_ sg13g2_buf_1
X_21175_ _02383_ _02360_ _02384_ VPWR VGND _01498_ sg13g2_mux2_1
X_21176_ \atbs_core_0.spike_memory_0.n2388_o[17]\ VPWR VGND _02385_ sg13g2_buf_1
X_21177_ _02385_ _02361_ _02384_ VPWR VGND _01499_ sg13g2_mux2_1
X_21178_ \atbs_core_0.spike_memory_0.n2388_o[18]\ VPWR VGND _02386_ sg13g2_buf_1
X_21179_ _02386_ _02364_ _02384_ VPWR VGND _01500_ sg13g2_mux2_1
X_21180_ \atbs_core_0.spike_memory_0.n2389_o[0]\ _02366_ _02384_ VPWR VGND _01501_ sg13g2_mux2_1
X_21181_ \atbs_core_0.spike_memory_0.n2361_o[1]\ _02232_ _02384_ VPWR VGND _01502_ sg13g2_mux2_1
X_21182_ \atbs_core_0.spike_memory_0.n2389_o[1]\ _02367_ _02384_ VPWR VGND _01503_ sg13g2_mux2_1
X_21183_ \atbs_core_0.spike_memory_0.n2389_o[2]\ _02368_ _02384_ VPWR VGND _01504_ sg13g2_mux2_1
X_21184_ \atbs_core_0.spike_memory_0.n2389_o[3]\ _02369_ _02384_ VPWR VGND _01505_ sg13g2_mux2_1
X_21185_ \atbs_core_0.spike_memory_0.n2389_o[4]\ _02370_ _02384_ VPWR VGND _01506_ sg13g2_mux2_1
X_21186_ \atbs_core_0.spike_memory_0.n2389_o[5]\ _02371_ _02384_ VPWR VGND _01507_ sg13g2_mux2_1
X_21187_ _02362_ VPWR VGND _02387_ sg13g2_buf_1
X_21188_ \atbs_core_0.spike_memory_0.n2389_o[6]\ _02372_ _02387_ VPWR VGND _01508_ sg13g2_mux2_1
X_21189_ \atbs_core_0.spike_memory_0.n2389_o[7]\ _02373_ _02387_ VPWR VGND _01509_ sg13g2_mux2_1
X_21190_ \atbs_core_0.spike_memory_0.n2389_o[8]\ _02375_ _02387_ VPWR VGND _01510_ sg13g2_mux2_1
X_21191_ \atbs_core_0.spike_memory_0.n2389_o[9]\ _02376_ _02387_ VPWR VGND _01511_ sg13g2_mux2_1
X_21192_ \atbs_core_0.spike_memory_0.n2389_o[10]\ _02377_ _02387_ VPWR VGND _01512_ sg13g2_mux2_1
X_21193_ \atbs_core_0.spike_memory_0.n2361_o[2]\ _02244_ _02387_ VPWR VGND _01513_ sg13g2_mux2_1
X_21194_ \atbs_core_0.spike_memory_0.n2358_o[5]\ \atbs_core_0.spike_memory_0.a_data[5]\ _02387_ VPWR VGND _01514_ sg13g2_mux2_1
X_21195_ \atbs_core_0.spike_memory_0.n2389_o[11]\ _02378_ _02387_ VPWR VGND _01515_ sg13g2_mux2_1
X_21196_ \atbs_core_0.spike_memory_0.n2389_o[12]\ _02379_ _02387_ VPWR VGND _01516_ sg13g2_mux2_1
X_21197_ \atbs_core_0.spike_memory_0.n2389_o[13]\ _02380_ _02387_ VPWR VGND _01517_ sg13g2_mux2_1
X_21198_ _02362_ VPWR VGND _02388_ sg13g2_buf_1
X_21199_ \atbs_core_0.spike_memory_0.n2389_o[14]\ _02381_ _02388_ VPWR VGND _01518_ sg13g2_mux2_1
X_21200_ \atbs_core_0.spike_memory_0.n2389_o[15]\ _02382_ _02388_ VPWR VGND _01519_ sg13g2_mux2_1
X_21201_ \atbs_core_0.spike_memory_0.n2389_o[16]\ _02383_ _02388_ VPWR VGND _01520_ sg13g2_mux2_1
X_21202_ \atbs_core_0.spike_memory_0.n2389_o[17]\ _02385_ _02388_ VPWR VGND _01521_ sg13g2_mux2_1
X_21203_ \atbs_core_0.spike_memory_0.n2389_o[18]\ _02386_ _02388_ VPWR VGND _01522_ sg13g2_mux2_1
X_21204_ \atbs_core_0.spike_memory_0.n2390_o[0]\ \atbs_core_0.spike_memory_0.n2389_o[0]\ _02388_ VPWR VGND _01523_ sg13g2_mux2_1
X_21205_ \atbs_core_0.spike_memory_0.n2390_o[1]\ \atbs_core_0.spike_memory_0.n2389_o[1]\ _02388_ VPWR VGND _01524_ sg13g2_mux2_1
X_21206_ \atbs_core_0.spike_memory_0.n2361_o[3]\ _02256_ _02388_ VPWR VGND _01525_ sg13g2_mux2_1
X_21207_ \atbs_core_0.spike_memory_0.n2390_o[2]\ \atbs_core_0.spike_memory_0.n2389_o[2]\ _02388_ VPWR VGND _01526_ sg13g2_mux2_1
X_21208_ \atbs_core_0.spike_memory_0.n2390_o[3]\ \atbs_core_0.spike_memory_0.n2389_o[3]\ _02388_ VPWR VGND _01527_ sg13g2_mux2_1
X_21209_ _02362_ VPWR VGND _02389_ sg13g2_buf_1
X_21210_ \atbs_core_0.spike_memory_0.n2390_o[4]\ \atbs_core_0.spike_memory_0.n2389_o[4]\ _02389_ VPWR VGND _01528_ sg13g2_mux2_1
X_21211_ \atbs_core_0.spike_memory_0.n2390_o[5]\ \atbs_core_0.spike_memory_0.n2389_o[5]\ _02389_ VPWR VGND _01529_ sg13g2_mux2_1
X_21212_ \atbs_core_0.spike_memory_0.n2390_o[6]\ \atbs_core_0.spike_memory_0.n2389_o[6]\ _02389_ VPWR VGND _01530_ sg13g2_mux2_1
X_21213_ \atbs_core_0.spike_memory_0.n2390_o[7]\ \atbs_core_0.spike_memory_0.n2389_o[7]\ _02389_ VPWR VGND _01531_ sg13g2_mux2_1
X_21214_ \atbs_core_0.spike_memory_0.n2390_o[8]\ \atbs_core_0.spike_memory_0.n2389_o[8]\ _02389_ VPWR VGND _01532_ sg13g2_mux2_1
X_21215_ \atbs_core_0.spike_memory_0.n2390_o[9]\ \atbs_core_0.spike_memory_0.n2389_o[9]\ _02389_ VPWR VGND _01533_ sg13g2_mux2_1
X_21216_ \atbs_core_0.spike_memory_0.n2390_o[10]\ \atbs_core_0.spike_memory_0.n2389_o[10]\ _02389_ VPWR VGND _01534_ sg13g2_mux2_1
X_21217_ \atbs_core_0.spike_memory_0.n2390_o[11]\ \atbs_core_0.spike_memory_0.n2389_o[11]\ _02389_ VPWR VGND _01535_ sg13g2_mux2_1
X_21218_ \atbs_core_0.spike_memory_0.n2361_o[4]\ _02268_ _02389_ VPWR VGND _01536_ sg13g2_mux2_1
X_21219_ \atbs_core_0.spike_memory_0.n2390_o[12]\ \atbs_core_0.spike_memory_0.n2389_o[12]\ _02389_ VPWR VGND _01537_ sg13g2_mux2_1
X_21220_ _02362_ VPWR VGND _02390_ sg13g2_buf_1
X_21221_ \atbs_core_0.spike_memory_0.n2390_o[13]\ \atbs_core_0.spike_memory_0.n2389_o[13]\ _02390_ VPWR VGND _01538_ sg13g2_mux2_1
X_21222_ \atbs_core_0.spike_memory_0.n2390_o[14]\ \atbs_core_0.spike_memory_0.n2389_o[14]\ _02390_ VPWR VGND _01539_ sg13g2_mux2_1
X_21223_ \atbs_core_0.spike_memory_0.n2390_o[15]\ \atbs_core_0.spike_memory_0.n2389_o[15]\ _02390_ VPWR VGND _01540_ sg13g2_mux2_1
X_21224_ \atbs_core_0.spike_memory_0.n2390_o[16]\ \atbs_core_0.spike_memory_0.n2389_o[16]\ _02390_ VPWR VGND _01541_ sg13g2_mux2_1
X_21225_ \atbs_core_0.spike_memory_0.n2390_o[17]\ \atbs_core_0.spike_memory_0.n2389_o[17]\ _02390_ VPWR VGND _01542_ sg13g2_mux2_1
X_21226_ \atbs_core_0.spike_memory_0.n2390_o[18]\ \atbs_core_0.spike_memory_0.n2389_o[18]\ _02390_ VPWR VGND _01543_ sg13g2_mux2_1
X_21227_ \atbs_core_0.spike_memory_0.n2391_o[0]\ VPWR VGND _02391_ sg13g2_buf_1
X_21228_ _02391_ \atbs_core_0.spike_memory_0.n2390_o[0]\ _02390_ VPWR VGND _01544_ sg13g2_mux2_1
X_21229_ \atbs_core_0.spike_memory_0.n2391_o[1]\ VPWR VGND _02392_ sg13g2_buf_1
X_21230_ _02392_ \atbs_core_0.spike_memory_0.n2390_o[1]\ _02390_ VPWR VGND _01545_ sg13g2_mux2_1
X_21231_ \atbs_core_0.spike_memory_0.n2391_o[2]\ \atbs_core_0.spike_memory_0.n2390_o[2]\ _02390_ VPWR VGND _01546_ sg13g2_mux2_1
X_21232_ \atbs_core_0.spike_memory_0.n2361_o[5]\ _02277_ _02390_ VPWR VGND _01547_ sg13g2_mux2_1
X_21233_ \atbs_core_0.spike_memory_0.n2391_o[3]\ VPWR VGND _02393_ sg13g2_buf_1
X_21234_ _02074_ VPWR VGND _02394_ sg13g2_buf_1
X_21235_ _02394_ VPWR VGND _02395_ sg13g2_buf_1
X_21236_ _02393_ \atbs_core_0.spike_memory_0.n2390_o[3]\ _02395_ VPWR VGND _01548_ sg13g2_mux2_1
X_21237_ \atbs_core_0.spike_memory_0.n2391_o[4]\ VPWR VGND _02396_ sg13g2_buf_1
X_21238_ _02396_ \atbs_core_0.spike_memory_0.n2390_o[4]\ _02395_ VPWR VGND _01549_ sg13g2_mux2_1
X_21239_ \atbs_core_0.spike_memory_0.n2391_o[5]\ \atbs_core_0.spike_memory_0.n2390_o[5]\ _02395_ VPWR VGND _01550_ sg13g2_mux2_1
X_21240_ \atbs_core_0.spike_memory_0.n2391_o[6]\ VPWR VGND _02397_ sg13g2_buf_1
X_21241_ _02397_ \atbs_core_0.spike_memory_0.n2390_o[6]\ _02395_ VPWR VGND _01551_ sg13g2_mux2_1
X_21242_ \atbs_core_0.spike_memory_0.n2391_o[7]\ VPWR VGND _02398_ sg13g2_buf_1
X_21243_ _02398_ \atbs_core_0.spike_memory_0.n2390_o[7]\ _02395_ VPWR VGND _01552_ sg13g2_mux2_1
X_21244_ \atbs_core_0.spike_memory_0.n2391_o[8]\ VPWR VGND _02399_ sg13g2_buf_1
X_21245_ _02399_ \atbs_core_0.spike_memory_0.n2390_o[8]\ _02395_ VPWR VGND _01553_ sg13g2_mux2_1
X_21246_ \atbs_core_0.spike_memory_0.n2391_o[9]\ VPWR VGND _02400_ sg13g2_buf_1
X_21247_ _02400_ \atbs_core_0.spike_memory_0.n2390_o[9]\ _02395_ VPWR VGND _01554_ sg13g2_mux2_1
X_21248_ \atbs_core_0.spike_memory_0.n2391_o[10]\ VPWR VGND _02401_ sg13g2_buf_1
X_21249_ _02401_ \atbs_core_0.spike_memory_0.n2390_o[10]\ _02395_ VPWR VGND _01555_ sg13g2_mux2_1
X_21250_ \atbs_core_0.spike_memory_0.n2391_o[11]\ VPWR VGND _02402_ sg13g2_buf_1
X_21251_ _02402_ \atbs_core_0.spike_memory_0.n2390_o[11]\ _02395_ VPWR VGND _01556_ sg13g2_mux2_1
X_21252_ \atbs_core_0.spike_memory_0.n2391_o[12]\ VPWR VGND _02403_ sg13g2_buf_1
X_21253_ _02403_ \atbs_core_0.spike_memory_0.n2390_o[12]\ _02395_ VPWR VGND _01557_ sg13g2_mux2_1
X_21254_ _02394_ VPWR VGND _02404_ sg13g2_buf_1
X_21255_ \atbs_core_0.spike_memory_0.n2361_o[6]\ _02280_ _02404_ VPWR VGND _01558_ sg13g2_mux2_1
X_21256_ \atbs_core_0.spike_memory_0.n2391_o[13]\ VPWR VGND _02405_ sg13g2_buf_1
X_21257_ _02405_ \atbs_core_0.spike_memory_0.n2390_o[13]\ _02404_ VPWR VGND _01559_ sg13g2_mux2_1
X_21258_ \atbs_core_0.spike_memory_0.n2391_o[14]\ VPWR VGND _02406_ sg13g2_buf_1
X_21259_ _02406_ \atbs_core_0.spike_memory_0.n2390_o[14]\ _02404_ VPWR VGND _01560_ sg13g2_mux2_1
X_21260_ \atbs_core_0.spike_memory_0.n2391_o[15]\ VPWR VGND _02407_ sg13g2_buf_1
X_21261_ _02407_ \atbs_core_0.spike_memory_0.n2390_o[15]\ _02404_ VPWR VGND _01561_ sg13g2_mux2_1
X_21262_ \atbs_core_0.spike_memory_0.n2391_o[16]\ VPWR VGND _02408_ sg13g2_buf_1
X_21263_ _02408_ \atbs_core_0.spike_memory_0.n2390_o[16]\ _02404_ VPWR VGND _01562_ sg13g2_mux2_1
X_21264_ \atbs_core_0.spike_memory_0.n2391_o[17]\ VPWR VGND _02409_ sg13g2_buf_1
X_21265_ _02409_ \atbs_core_0.spike_memory_0.n2390_o[17]\ _02404_ VPWR VGND _01563_ sg13g2_mux2_1
X_21266_ \atbs_core_0.spike_memory_0.n2391_o[18]\ VPWR VGND _02410_ sg13g2_buf_1
X_21267_ _02410_ \atbs_core_0.spike_memory_0.n2390_o[18]\ _02404_ VPWR VGND _01564_ sg13g2_mux2_1
X_21268_ \atbs_core_0.spike_memory_0.n2392_o[0]\ VPWR VGND _02411_ sg13g2_buf_1
X_21269_ _02411_ _02391_ _02404_ VPWR VGND _01565_ sg13g2_mux2_1
X_21270_ \atbs_core_0.spike_memory_0.n2392_o[1]\ VPWR VGND _02412_ sg13g2_buf_1
X_21271_ _02412_ _02392_ _02404_ VPWR VGND _01566_ sg13g2_mux2_1
X_21272_ \atbs_core_0.spike_memory_0.n2392_o[2]\ \atbs_core_0.spike_memory_0.n2391_o[2]\ _02404_ VPWR VGND _01567_ sg13g2_mux2_1
X_21273_ \atbs_core_0.spike_memory_0.n2392_o[3]\ VPWR VGND _02413_ sg13g2_buf_1
X_21274_ _02394_ VPWR VGND _02414_ sg13g2_buf_1
X_21275_ _02413_ _02393_ _02414_ VPWR VGND _01568_ sg13g2_mux2_1
X_21276_ \atbs_core_0.spike_memory_0.n2361_o[7]\ _02282_ _02414_ VPWR VGND _01569_ sg13g2_mux2_1
X_21277_ \atbs_core_0.spike_memory_0.n2392_o[4]\ VPWR VGND _02415_ sg13g2_buf_1
X_21278_ _02415_ _02396_ _02414_ VPWR VGND _01570_ sg13g2_mux2_1
X_21279_ \atbs_core_0.spike_memory_0.n2392_o[5]\ \atbs_core_0.spike_memory_0.n2391_o[5]\ _02414_ VPWR VGND _01571_ sg13g2_mux2_1
X_21280_ \atbs_core_0.spike_memory_0.n2392_o[6]\ VPWR VGND _02416_ sg13g2_buf_1
X_21281_ _02416_ _02397_ _02414_ VPWR VGND _01572_ sg13g2_mux2_1
X_21282_ \atbs_core_0.spike_memory_0.n2392_o[7]\ VPWR VGND _02417_ sg13g2_buf_1
X_21283_ _02417_ _02398_ _02414_ VPWR VGND _01573_ sg13g2_mux2_1
X_21284_ \atbs_core_0.spike_memory_0.n2392_o[8]\ VPWR VGND _02418_ sg13g2_buf_1
X_21285_ _02418_ _02399_ _02414_ VPWR VGND _01574_ sg13g2_mux2_1
X_21286_ \atbs_core_0.spike_memory_0.n2392_o[9]\ VPWR VGND _02419_ sg13g2_buf_1
X_21287_ _02419_ _02400_ _02414_ VPWR VGND _01575_ sg13g2_mux2_1
X_21288_ \atbs_core_0.spike_memory_0.n2392_o[10]\ VPWR VGND _02420_ sg13g2_buf_1
X_21289_ _02420_ _02401_ _02414_ VPWR VGND _01576_ sg13g2_mux2_1
X_21290_ \atbs_core_0.spike_memory_0.n2392_o[11]\ VPWR VGND _02421_ sg13g2_buf_1
X_21291_ _02421_ _02402_ _02414_ VPWR VGND _01577_ sg13g2_mux2_1
X_21292_ \atbs_core_0.spike_memory_0.n2392_o[12]\ VPWR VGND _02422_ sg13g2_buf_1
X_21293_ _02394_ VPWR VGND _02423_ sg13g2_buf_1
X_21294_ _02422_ _02403_ _02423_ VPWR VGND _01578_ sg13g2_mux2_1
X_21295_ \atbs_core_0.spike_memory_0.n2392_o[13]\ VPWR VGND _02424_ sg13g2_buf_1
X_21296_ _02424_ _02405_ _02423_ VPWR VGND _01579_ sg13g2_mux2_1
X_21297_ \atbs_core_0.spike_memory_0.n2361_o[8]\ _02285_ _02423_ VPWR VGND _01580_ sg13g2_mux2_1
X_21298_ \atbs_core_0.spike_memory_0.n2392_o[14]\ VPWR VGND _02425_ sg13g2_buf_1
X_21299_ _02425_ _02406_ _02423_ VPWR VGND _01581_ sg13g2_mux2_1
X_21300_ \atbs_core_0.spike_memory_0.n2392_o[15]\ VPWR VGND _02426_ sg13g2_buf_1
X_21301_ _02426_ _02407_ _02423_ VPWR VGND _01582_ sg13g2_mux2_1
X_21302_ \atbs_core_0.spike_memory_0.n2392_o[16]\ VPWR VGND _02427_ sg13g2_buf_1
X_21303_ _02427_ _02408_ _02423_ VPWR VGND _01583_ sg13g2_mux2_1
X_21304_ \atbs_core_0.spike_memory_0.n2392_o[17]\ VPWR VGND _02428_ sg13g2_buf_1
X_21305_ _02428_ _02409_ _02423_ VPWR VGND _01584_ sg13g2_mux2_1
X_21306_ \atbs_core_0.spike_memory_0.n2392_o[18]\ VPWR VGND _02429_ sg13g2_buf_1
X_21307_ _02429_ _02410_ _02423_ VPWR VGND _01585_ sg13g2_mux2_1
X_21308_ \atbs_core_0.spike_memory_0.n2393_o[0]\ VPWR VGND _02430_ sg13g2_inv_1
X_21309_ _02411_ _02217_ VPWR VGND _02431_ sg13g2_nand2_1
X_21310_ _02430_ _02208_ _02431_ VPWR VGND _01586_ sg13g2_o21ai_1
X_21311_ \atbs_core_0.spike_memory_0.n2393_o[1]\ VPWR VGND _02432_ sg13g2_inv_1
X_21312_ _12513_ VPWR VGND _02433_ sg13g2_buf_1
X_21313_ _02412_ _02217_ VPWR VGND _02434_ sg13g2_nand2_1
X_21314_ _02432_ _02433_ _02434_ VPWR VGND _01587_ sg13g2_o21ai_1
X_21315_ \atbs_core_0.spike_memory_0.n2393_o[2]\ VPWR VGND _02435_ sg13g2_inv_1
X_21316_ \atbs_core_0.spike_memory_0.n2392_o[2]\ _02217_ VPWR VGND _02436_ sg13g2_nand2_1
X_21317_ _02435_ _02433_ _02436_ VPWR VGND _01588_ sg13g2_o21ai_1
X_21318_ \atbs_core_0.spike_memory_0.n2393_o[3]\ VPWR VGND _02437_ sg13g2_inv_1
X_21319_ _02413_ _02217_ VPWR VGND _02438_ sg13g2_nand2_1
X_21320_ _02437_ _02433_ _02438_ VPWR VGND _01589_ sg13g2_o21ai_1
X_21321_ \atbs_core_0.spike_memory_0.n2393_o[4]\ VPWR VGND _02439_ sg13g2_inv_1
X_21322_ _02415_ _02217_ VPWR VGND _02440_ sg13g2_nand2_1
X_21323_ _02439_ _02433_ _02440_ VPWR VGND _01590_ sg13g2_o21ai_1
X_21324_ \atbs_core_0.spike_memory_0.n2361_o[9]\ _02292_ _02423_ VPWR VGND _01591_ sg13g2_mux2_1
X_21325_ \atbs_core_0.spike_memory_0.n2393_o[5]\ VPWR VGND _02441_ sg13g2_inv_1
X_21326_ _02191_ VPWR VGND _02442_ sg13g2_buf_1
X_21327_ \atbs_core_0.spike_memory_0.n2392_o[5]\ _02442_ VPWR VGND _02443_ sg13g2_nand2_1
X_21328_ _02441_ _02433_ _02443_ VPWR VGND _01592_ sg13g2_o21ai_1
X_21329_ \atbs_core_0.spike_memory_0.n2393_o[6]\ VPWR VGND _02444_ sg13g2_inv_1
X_21330_ _02416_ _02442_ VPWR VGND _02445_ sg13g2_nand2_1
X_21331_ _02444_ _02433_ _02445_ VPWR VGND _01593_ sg13g2_o21ai_1
X_21332_ \atbs_core_0.spike_memory_0.n2393_o[7]\ VPWR VGND _02446_ sg13g2_inv_1
X_21333_ _02417_ _02442_ VPWR VGND _02447_ sg13g2_nand2_1
X_21334_ _02446_ _02433_ _02447_ VPWR VGND _01594_ sg13g2_o21ai_1
X_21335_ \atbs_core_0.spike_memory_0.n2393_o[8]\ VPWR VGND _02448_ sg13g2_inv_1
X_21336_ _02418_ _02442_ VPWR VGND _02449_ sg13g2_nand2_1
X_21337_ _02448_ _02433_ _02449_ VPWR VGND _01595_ sg13g2_o21ai_1
X_21338_ \atbs_core_0.spike_memory_0.n2393_o[9]\ VPWR VGND _02450_ sg13g2_inv_1
X_21339_ _02419_ _02442_ VPWR VGND _02451_ sg13g2_nand2_1
X_21340_ _02450_ _02433_ _02451_ VPWR VGND _01596_ sg13g2_o21ai_1
X_21341_ \atbs_core_0.spike_memory_0.n2393_o[10]\ VPWR VGND _02452_ sg13g2_inv_1
X_21342_ _02420_ _02442_ VPWR VGND _02453_ sg13g2_nand2_1
X_21343_ _02452_ _02433_ _02453_ VPWR VGND _01597_ sg13g2_o21ai_1
X_21344_ \atbs_core_0.spike_memory_0.n2393_o[11]\ VPWR VGND _02454_ sg13g2_inv_1
X_21345_ _12513_ VPWR VGND _02455_ sg13g2_buf_1
X_21346_ _02421_ _02442_ VPWR VGND _02456_ sg13g2_nand2_1
X_21347_ _02454_ _02455_ _02456_ VPWR VGND _01598_ sg13g2_o21ai_1
X_21348_ \atbs_core_0.spike_memory_0.n2393_o[12]\ VPWR VGND _02457_ sg13g2_inv_1
X_21349_ _02422_ _02442_ VPWR VGND _02458_ sg13g2_nand2_1
X_21350_ _02457_ _02455_ _02458_ VPWR VGND _01599_ sg13g2_o21ai_1
X_21351_ \atbs_core_0.spike_memory_0.n2393_o[13]\ VPWR VGND _02459_ sg13g2_inv_1
X_21352_ _02424_ _02442_ VPWR VGND _02460_ sg13g2_nand2_1
X_21353_ _02459_ _02455_ _02460_ VPWR VGND _01600_ sg13g2_o21ai_1
X_21354_ \atbs_core_0.spike_memory_0.n2393_o[14]\ VPWR VGND _02461_ sg13g2_inv_1
X_21355_ _02425_ _02442_ VPWR VGND _02462_ sg13g2_nand2_1
X_21356_ _02461_ _02455_ _02462_ VPWR VGND _01601_ sg13g2_o21ai_1
X_21357_ \atbs_core_0.spike_memory_0.n2361_o[10]\ _02304_ _02423_ VPWR VGND _01602_ sg13g2_mux2_1
X_21358_ \atbs_core_0.spike_memory_0.n2393_o[15]\ VPWR VGND _02463_ sg13g2_inv_1
X_21359_ _02191_ VPWR VGND _02464_ sg13g2_buf_1
X_21360_ _02426_ _02464_ VPWR VGND _02465_ sg13g2_nand2_1
X_21361_ _02463_ _02455_ _02465_ VPWR VGND _01603_ sg13g2_o21ai_1
X_21362_ \atbs_core_0.spike_memory_0.n2393_o[16]\ VPWR VGND _02466_ sg13g2_inv_1
X_21363_ _02427_ _02464_ VPWR VGND _02467_ sg13g2_nand2_1
X_21364_ _02466_ _02455_ _02467_ VPWR VGND _01604_ sg13g2_o21ai_1
X_21365_ \atbs_core_0.spike_memory_0.n2393_o[17]\ VPWR VGND _02468_ sg13g2_inv_1
X_21366_ _02428_ _02464_ VPWR VGND _02469_ sg13g2_nand2_1
X_21367_ _02468_ _02455_ _02469_ VPWR VGND _01605_ sg13g2_o21ai_1
X_21368_ \atbs_core_0.spike_memory_0.n2393_o[18]\ VPWR VGND _02470_ sg13g2_inv_1
X_21369_ _02429_ _02464_ VPWR VGND _02471_ sg13g2_nand2_1
X_21370_ _02470_ _02455_ _02471_ VPWR VGND _01606_ sg13g2_o21ai_1
X_21371_ _02394_ VPWR VGND _02472_ sg13g2_buf_1
X_21372_ \atbs_core_0.spike_memory_0.n2394_o[0]\ \atbs_core_0.spike_memory_0.n2393_o[0]\ _02472_ VPWR VGND _01607_ sg13g2_mux2_1
X_21373_ \atbs_core_0.spike_memory_0.n2394_o[1]\ \atbs_core_0.spike_memory_0.n2393_o[1]\ _02472_ VPWR VGND _01608_ sg13g2_mux2_1
X_21374_ \atbs_core_0.spike_memory_0.n2394_o[2]\ \atbs_core_0.spike_memory_0.n2393_o[2]\ _02472_ VPWR VGND _01609_ sg13g2_mux2_1
X_21375_ \atbs_core_0.spike_memory_0.n2394_o[3]\ \atbs_core_0.spike_memory_0.n2393_o[3]\ _02472_ VPWR VGND _01610_ sg13g2_mux2_1
X_21376_ \atbs_core_0.spike_memory_0.n2394_o[4]\ \atbs_core_0.spike_memory_0.n2393_o[4]\ _02472_ VPWR VGND _01611_ sg13g2_mux2_1
X_21377_ \atbs_core_0.spike_memory_0.n2394_o[5]\ \atbs_core_0.spike_memory_0.n2393_o[5]\ _02472_ VPWR VGND _01612_ sg13g2_mux2_1
X_21378_ \atbs_core_0.spike_memory_0.n2361_o[11]\ _02316_ _02472_ VPWR VGND _01613_ sg13g2_mux2_1
X_21379_ \atbs_core_0.spike_memory_0.n2394_o[6]\ \atbs_core_0.spike_memory_0.n2393_o[6]\ _02472_ VPWR VGND _01614_ sg13g2_mux2_1
X_21380_ \atbs_core_0.spike_memory_0.n2394_o[7]\ \atbs_core_0.spike_memory_0.n2393_o[7]\ _02472_ VPWR VGND _01615_ sg13g2_mux2_1
X_21381_ \atbs_core_0.spike_memory_0.n2394_o[8]\ \atbs_core_0.spike_memory_0.n2393_o[8]\ _02472_ VPWR VGND _01616_ sg13g2_mux2_1
X_21382_ _02394_ VPWR VGND _02473_ sg13g2_buf_1
X_21383_ \atbs_core_0.spike_memory_0.n2394_o[9]\ \atbs_core_0.spike_memory_0.n2393_o[9]\ _02473_ VPWR VGND _01617_ sg13g2_mux2_1
X_21384_ \atbs_core_0.spike_memory_0.n2394_o[10]\ \atbs_core_0.spike_memory_0.n2393_o[10]\ _02473_ VPWR VGND _01618_ sg13g2_mux2_1
X_21385_ \atbs_core_0.spike_memory_0.n2394_o[11]\ \atbs_core_0.spike_memory_0.n2393_o[11]\ _02473_ VPWR VGND _01619_ sg13g2_mux2_1
X_21386_ \atbs_core_0.spike_memory_0.n2394_o[12]\ \atbs_core_0.spike_memory_0.n2393_o[12]\ _02473_ VPWR VGND _01620_ sg13g2_mux2_1
X_21387_ \atbs_core_0.spike_memory_0.n2394_o[13]\ \atbs_core_0.spike_memory_0.n2393_o[13]\ _02473_ VPWR VGND _01621_ sg13g2_mux2_1
X_21388_ \atbs_core_0.spike_memory_0.n2394_o[14]\ \atbs_core_0.spike_memory_0.n2393_o[14]\ _02473_ VPWR VGND _01622_ sg13g2_mux2_1
X_21389_ \atbs_core_0.spike_memory_0.n2394_o[15]\ \atbs_core_0.spike_memory_0.n2393_o[15]\ _02473_ VPWR VGND _01623_ sg13g2_mux2_1
X_21390_ \atbs_core_0.spike_memory_0.n2361_o[12]\ _02329_ _02473_ VPWR VGND _01624_ sg13g2_mux2_1
X_21391_ \atbs_core_0.spike_memory_0.n2358_o[6]\ \atbs_core_0.spike_memory_0.a_data[6]\ _02473_ VPWR VGND _01625_ sg13g2_mux2_1
X_21392_ \atbs_core_0.spike_memory_0.n2394_o[16]\ \atbs_core_0.spike_memory_0.n2393_o[16]\ _02473_ VPWR VGND _01626_ sg13g2_mux2_1
X_21393_ _02394_ VPWR VGND _02474_ sg13g2_buf_1
X_21394_ \atbs_core_0.spike_memory_0.n2394_o[17]\ \atbs_core_0.spike_memory_0.n2393_o[17]\ _02474_ VPWR VGND _01627_ sg13g2_mux2_1
X_21395_ \atbs_core_0.spike_memory_0.n2394_o[18]\ \atbs_core_0.spike_memory_0.n2393_o[18]\ _02474_ VPWR VGND _01628_ sg13g2_mux2_1
X_21396_ \atbs_core_0.spike_memory_0.n2395_o[0]\ VPWR VGND _02475_ sg13g2_buf_1
X_21397_ _02475_ \atbs_core_0.spike_memory_0.n2394_o[0]\ _02474_ VPWR VGND _01629_ sg13g2_mux2_1
X_21398_ \atbs_core_0.spike_memory_0.n2395_o[1]\ VPWR VGND _02476_ sg13g2_buf_1
X_21399_ _02476_ \atbs_core_0.spike_memory_0.n2394_o[1]\ _02474_ VPWR VGND _01630_ sg13g2_mux2_1
X_21400_ \atbs_core_0.spike_memory_0.n2395_o[2]\ VPWR VGND _02477_ sg13g2_buf_1
X_21401_ _02477_ \atbs_core_0.spike_memory_0.n2394_o[2]\ _02474_ VPWR VGND _01631_ sg13g2_mux2_1
X_21402_ \atbs_core_0.spike_memory_0.n2395_o[3]\ VPWR VGND _02478_ sg13g2_buf_1
X_21403_ _02478_ \atbs_core_0.spike_memory_0.n2394_o[3]\ _02474_ VPWR VGND _01632_ sg13g2_mux2_1
X_21404_ \atbs_core_0.spike_memory_0.n2395_o[4]\ VPWR VGND _02479_ sg13g2_buf_1
X_21405_ _02479_ \atbs_core_0.spike_memory_0.n2394_o[4]\ _02474_ VPWR VGND _01633_ sg13g2_mux2_1
X_21406_ \atbs_core_0.spike_memory_0.n2395_o[5]\ VPWR VGND _02480_ sg13g2_buf_1
X_21407_ _02480_ \atbs_core_0.spike_memory_0.n2394_o[5]\ _02474_ VPWR VGND _01634_ sg13g2_mux2_1
X_21408_ \atbs_core_0.spike_memory_0.n2395_o[6]\ VPWR VGND _02481_ sg13g2_buf_1
X_21409_ _02481_ \atbs_core_0.spike_memory_0.n2394_o[6]\ _02474_ VPWR VGND _01635_ sg13g2_mux2_1
X_21410_ \atbs_core_0.spike_memory_0.n2361_o[13]\ _02334_ _02474_ VPWR VGND _01636_ sg13g2_mux2_1
X_21411_ \atbs_core_0.spike_memory_0.n2395_o[7]\ VPWR VGND _02482_ sg13g2_buf_1
X_21412_ _12511_ VPWR VGND _02483_ sg13g2_buf_1
X_21413_ _02483_ VPWR VGND _02484_ sg13g2_buf_1
X_21414_ _02482_ \atbs_core_0.spike_memory_0.n2394_o[7]\ _02484_ VPWR VGND _01637_ sg13g2_mux2_1
X_21415_ \atbs_core_0.spike_memory_0.n2395_o[8]\ VPWR VGND _02485_ sg13g2_buf_1
X_21416_ _02485_ \atbs_core_0.spike_memory_0.n2394_o[8]\ _02484_ VPWR VGND _01638_ sg13g2_mux2_1
X_21417_ \atbs_core_0.spike_memory_0.n2395_o[9]\ VPWR VGND _02486_ sg13g2_buf_1
X_21418_ _02486_ \atbs_core_0.spike_memory_0.n2394_o[9]\ _02484_ VPWR VGND _01639_ sg13g2_mux2_1
X_21419_ \atbs_core_0.spike_memory_0.n2395_o[10]\ VPWR VGND _02487_ sg13g2_buf_1
X_21420_ _02487_ \atbs_core_0.spike_memory_0.n2394_o[10]\ _02484_ VPWR VGND _01640_ sg13g2_mux2_1
X_21421_ \atbs_core_0.spike_memory_0.n2395_o[11]\ VPWR VGND _02488_ sg13g2_buf_1
X_21422_ _02488_ \atbs_core_0.spike_memory_0.n2394_o[11]\ _02484_ VPWR VGND _01641_ sg13g2_mux2_1
X_21423_ \atbs_core_0.spike_memory_0.n2395_o[12]\ VPWR VGND _02489_ sg13g2_buf_1
X_21424_ _02489_ \atbs_core_0.spike_memory_0.n2394_o[12]\ _02484_ VPWR VGND _01642_ sg13g2_mux2_1
X_21425_ \atbs_core_0.spike_memory_0.n2395_o[13]\ VPWR VGND _02490_ sg13g2_buf_1
X_21426_ _02490_ \atbs_core_0.spike_memory_0.n2394_o[13]\ _02484_ VPWR VGND _01643_ sg13g2_mux2_1
X_21427_ \atbs_core_0.spike_memory_0.n2395_o[14]\ VPWR VGND _02491_ sg13g2_buf_1
X_21428_ _02491_ \atbs_core_0.spike_memory_0.n2394_o[14]\ _02484_ VPWR VGND _01644_ sg13g2_mux2_1
X_21429_ \atbs_core_0.spike_memory_0.n2395_o[15]\ VPWR VGND _02492_ sg13g2_buf_1
X_21430_ _02492_ \atbs_core_0.spike_memory_0.n2394_o[15]\ _02484_ VPWR VGND _01645_ sg13g2_mux2_1
X_21431_ \atbs_core_0.spike_memory_0.n2395_o[16]\ VPWR VGND _02493_ sg13g2_buf_1
X_21432_ _02493_ \atbs_core_0.spike_memory_0.n2394_o[16]\ _02484_ VPWR VGND _01646_ sg13g2_mux2_1
X_21433_ _02483_ VPWR VGND _02494_ sg13g2_buf_1
X_21434_ \atbs_core_0.spike_memory_0.n2361_o[14]\ _02336_ _02494_ VPWR VGND _01647_ sg13g2_mux2_1
X_21435_ \atbs_core_0.spike_memory_0.n2395_o[17]\ VPWR VGND _02495_ sg13g2_buf_1
X_21436_ _02495_ \atbs_core_0.spike_memory_0.n2394_o[17]\ _02494_ VPWR VGND _01648_ sg13g2_mux2_1
X_21437_ \atbs_core_0.spike_memory_0.n2395_o[18]\ VPWR VGND _02496_ sg13g2_buf_1
X_21438_ _02496_ \atbs_core_0.spike_memory_0.n2394_o[18]\ _02494_ VPWR VGND _01649_ sg13g2_mux2_1
X_21439_ \atbs_core_0.spike_memory_0.n2396_o[0]\ VPWR VGND _02497_ sg13g2_buf_1
X_21440_ _02497_ _02475_ _02494_ VPWR VGND _01650_ sg13g2_mux2_1
X_21441_ \atbs_core_0.spike_memory_0.n2396_o[1]\ VPWR VGND _02498_ sg13g2_buf_1
X_21442_ _02498_ _02476_ _02494_ VPWR VGND _01651_ sg13g2_mux2_1
X_21443_ \atbs_core_0.spike_memory_0.n2396_o[2]\ VPWR VGND _02499_ sg13g2_buf_1
X_21444_ _02499_ _02477_ _02494_ VPWR VGND _01652_ sg13g2_mux2_1
X_21445_ \atbs_core_0.spike_memory_0.n2396_o[3]\ VPWR VGND _02500_ sg13g2_buf_1
X_21446_ _02500_ _02478_ _02494_ VPWR VGND _01653_ sg13g2_mux2_1
X_21447_ \atbs_core_0.spike_memory_0.n2396_o[4]\ VPWR VGND _02501_ sg13g2_buf_1
X_21448_ _02501_ _02479_ _02494_ VPWR VGND _01654_ sg13g2_mux2_1
X_21449_ \atbs_core_0.spike_memory_0.n2396_o[5]\ VPWR VGND _02502_ sg13g2_buf_1
X_21450_ _02502_ _02480_ _02494_ VPWR VGND _01655_ sg13g2_mux2_1
X_21451_ \atbs_core_0.spike_memory_0.n2396_o[6]\ VPWR VGND _02503_ sg13g2_buf_1
X_21452_ _02503_ _02481_ _02494_ VPWR VGND _01656_ sg13g2_mux2_1
X_21453_ \atbs_core_0.spike_memory_0.n2396_o[7]\ VPWR VGND _02504_ sg13g2_buf_1
X_21454_ _02483_ VPWR VGND _02505_ sg13g2_buf_1
X_21455_ _02504_ _02482_ _02505_ VPWR VGND _01657_ sg13g2_mux2_1
X_21456_ \atbs_core_0.spike_memory_0.n2361_o[15]\ _02338_ _02505_ VPWR VGND _01658_ sg13g2_mux2_1
X_21457_ \atbs_core_0.spike_memory_0.n2396_o[8]\ VPWR VGND _02506_ sg13g2_buf_1
X_21458_ _02506_ _02485_ _02505_ VPWR VGND _01659_ sg13g2_mux2_1
X_21459_ \atbs_core_0.spike_memory_0.n2396_o[9]\ VPWR VGND _02507_ sg13g2_buf_1
X_21460_ _02507_ _02486_ _02505_ VPWR VGND _01660_ sg13g2_mux2_1
X_21461_ \atbs_core_0.spike_memory_0.n2396_o[10]\ VPWR VGND _02508_ sg13g2_buf_1
X_21462_ _02508_ _02487_ _02505_ VPWR VGND _01661_ sg13g2_mux2_1
X_21463_ \atbs_core_0.spike_memory_0.n2396_o[11]\ VPWR VGND _02509_ sg13g2_buf_1
X_21464_ _02509_ _02488_ _02505_ VPWR VGND _01662_ sg13g2_mux2_1
X_21465_ \atbs_core_0.spike_memory_0.n2396_o[12]\ VPWR VGND _02510_ sg13g2_buf_1
X_21466_ _02510_ _02489_ _02505_ VPWR VGND _01663_ sg13g2_mux2_1
X_21467_ \atbs_core_0.spike_memory_0.n2396_o[13]\ VPWR VGND _02511_ sg13g2_buf_1
X_21468_ _02511_ _02490_ _02505_ VPWR VGND _01664_ sg13g2_mux2_1
X_21469_ \atbs_core_0.spike_memory_0.n2396_o[14]\ VPWR VGND _02512_ sg13g2_buf_1
X_21470_ _02512_ _02491_ _02505_ VPWR VGND _01665_ sg13g2_mux2_1
X_21471_ \atbs_core_0.spike_memory_0.n2396_o[15]\ VPWR VGND _02513_ sg13g2_buf_1
X_21472_ _02513_ _02492_ _02505_ VPWR VGND _01666_ sg13g2_mux2_1
X_21473_ \atbs_core_0.spike_memory_0.n2396_o[16]\ VPWR VGND _02514_ sg13g2_buf_1
X_21474_ _02483_ VPWR VGND _02515_ sg13g2_buf_1
X_21475_ _02514_ _02493_ _02515_ VPWR VGND _01667_ sg13g2_mux2_1
X_21476_ \atbs_core_0.spike_memory_0.n2396_o[17]\ VPWR VGND _02516_ sg13g2_buf_1
X_21477_ _02516_ _02495_ _02515_ VPWR VGND _01668_ sg13g2_mux2_1
X_21478_ \atbs_core_0.spike_memory_0.n2361_o[16]\ _02340_ _02515_ VPWR VGND _01669_ sg13g2_mux2_1
X_21479_ \atbs_core_0.spike_memory_0.n2396_o[18]\ VPWR VGND _02517_ sg13g2_buf_1
X_21480_ _02517_ _02496_ _02515_ VPWR VGND _01670_ sg13g2_mux2_1
X_21481_ \atbs_core_0.spike_memory_0.n2397_o[0]\ _02497_ _02515_ VPWR VGND _01671_ sg13g2_mux2_1
X_21482_ \atbs_core_0.spike_memory_0.n2397_o[1]\ _02498_ _02515_ VPWR VGND _01672_ sg13g2_mux2_1
X_21483_ \atbs_core_0.spike_memory_0.n2397_o[2]\ _02499_ _02515_ VPWR VGND _01673_ sg13g2_mux2_1
X_21484_ \atbs_core_0.spike_memory_0.n2397_o[3]\ _02500_ _02515_ VPWR VGND _01674_ sg13g2_mux2_1
X_21485_ \atbs_core_0.spike_memory_0.n2397_o[4]\ _02501_ _02515_ VPWR VGND _01675_ sg13g2_mux2_1
X_21486_ \atbs_core_0.spike_memory_0.n2397_o[5]\ _02502_ _02515_ VPWR VGND _01676_ sg13g2_mux2_1
X_21487_ _02483_ VPWR VGND _02518_ sg13g2_buf_1
X_21488_ \atbs_core_0.spike_memory_0.n2397_o[6]\ _02503_ _02518_ VPWR VGND _01677_ sg13g2_mux2_1
X_21489_ \atbs_core_0.spike_memory_0.n2397_o[7]\ _02504_ _02518_ VPWR VGND _01678_ sg13g2_mux2_1
X_21490_ \atbs_core_0.spike_memory_0.n2397_o[8]\ _02506_ _02518_ VPWR VGND _01679_ sg13g2_mux2_1
X_21491_ \atbs_core_0.spike_memory_0.n2361_o[17]\ _02352_ _02518_ VPWR VGND _01680_ sg13g2_mux2_1
X_21492_ \atbs_core_0.spike_memory_0.n2397_o[9]\ _02507_ _02518_ VPWR VGND _01681_ sg13g2_mux2_1
X_21493_ \atbs_core_0.spike_memory_0.n2397_o[10]\ _02508_ _02518_ VPWR VGND _01682_ sg13g2_mux2_1
X_21494_ \atbs_core_0.spike_memory_0.n2397_o[11]\ _02509_ _02518_ VPWR VGND _01683_ sg13g2_mux2_1
X_21495_ \atbs_core_0.spike_memory_0.n2397_o[12]\ _02510_ _02518_ VPWR VGND _01684_ sg13g2_mux2_1
X_21496_ \atbs_core_0.spike_memory_0.n2397_o[13]\ _02511_ _02518_ VPWR VGND _01685_ sg13g2_mux2_1
X_21497_ \atbs_core_0.spike_memory_0.n2397_o[14]\ _02512_ _02518_ VPWR VGND _01686_ sg13g2_mux2_1
X_21498_ _02483_ VPWR VGND _02519_ sg13g2_buf_1
X_21499_ \atbs_core_0.spike_memory_0.n2397_o[15]\ _02513_ _02519_ VPWR VGND _01687_ sg13g2_mux2_1
X_21500_ \atbs_core_0.spike_memory_0.n2397_o[16]\ _02514_ _02519_ VPWR VGND _01688_ sg13g2_mux2_1
X_21501_ \atbs_core_0.spike_memory_0.n2397_o[17]\ _02516_ _02519_ VPWR VGND _01689_ sg13g2_mux2_1
X_21502_ \atbs_core_0.spike_memory_0.n2397_o[18]\ _02517_ _02519_ VPWR VGND _01690_ sg13g2_mux2_1
X_21503_ \atbs_core_0.spike_memory_0.n2361_o[18]\ _02365_ _02519_ VPWR VGND _01691_ sg13g2_mux2_1
X_21504_ \atbs_core_0.spike_memory_0.n2398_o[0]\ \atbs_core_0.spike_memory_0.n2397_o[0]\ _02519_ VPWR VGND _01692_ sg13g2_mux2_1
X_21505_ \atbs_core_0.spike_memory_0.n2398_o[1]\ \atbs_core_0.spike_memory_0.n2397_o[1]\ _02519_ VPWR VGND _01693_ sg13g2_mux2_1
X_21506_ \atbs_core_0.spike_memory_0.n2398_o[2]\ \atbs_core_0.spike_memory_0.n2397_o[2]\ _02519_ VPWR VGND _01694_ sg13g2_mux2_1
X_21507_ \atbs_core_0.spike_memory_0.n2398_o[3]\ \atbs_core_0.spike_memory_0.n2397_o[3]\ _02519_ VPWR VGND _01695_ sg13g2_mux2_1
X_21508_ \atbs_core_0.spike_memory_0.n2398_o[4]\ \atbs_core_0.spike_memory_0.n2397_o[4]\ _02519_ VPWR VGND _01696_ sg13g2_mux2_1
X_21509_ _02483_ VPWR VGND _02520_ sg13g2_buf_1
X_21510_ \atbs_core_0.spike_memory_0.n2398_o[5]\ \atbs_core_0.spike_memory_0.n2397_o[5]\ _02520_ VPWR VGND _01697_ sg13g2_mux2_1
X_21511_ \atbs_core_0.spike_memory_0.n2398_o[6]\ \atbs_core_0.spike_memory_0.n2397_o[6]\ _02520_ VPWR VGND _01698_ sg13g2_mux2_1
X_21512_ \atbs_core_0.spike_memory_0.n2398_o[7]\ \atbs_core_0.spike_memory_0.n2397_o[7]\ _02520_ VPWR VGND _01699_ sg13g2_mux2_1
X_21513_ \atbs_core_0.spike_memory_0.n2398_o[8]\ \atbs_core_0.spike_memory_0.n2397_o[8]\ _02520_ VPWR VGND _01700_ sg13g2_mux2_1
X_21514_ \atbs_core_0.spike_memory_0.n2398_o[9]\ \atbs_core_0.spike_memory_0.n2397_o[9]\ _02520_ VPWR VGND _01701_ sg13g2_mux2_1
X_21515_ \atbs_core_0.spike_memory_0.n2362_o[0]\ \atbs_core_0.spike_memory_0.n2361_o[0]\ _02520_ VPWR VGND _01702_ sg13g2_mux2_1
X_21516_ \atbs_core_0.spike_memory_0.n2398_o[10]\ \atbs_core_0.spike_memory_0.n2397_o[10]\ _02520_ VPWR VGND _01703_ sg13g2_mux2_1
X_21517_ \atbs_core_0.spike_memory_0.n2398_o[11]\ \atbs_core_0.spike_memory_0.n2397_o[11]\ _02520_ VPWR VGND _01704_ sg13g2_mux2_1
X_21518_ \atbs_core_0.spike_memory_0.n2398_o[12]\ \atbs_core_0.spike_memory_0.n2397_o[12]\ _02520_ VPWR VGND _01705_ sg13g2_mux2_1
X_21519_ \atbs_core_0.spike_memory_0.n2398_o[13]\ \atbs_core_0.spike_memory_0.n2397_o[13]\ _02520_ VPWR VGND _01706_ sg13g2_mux2_1
X_21520_ _12511_ VPWR VGND _02521_ sg13g2_buf_1
X_21521_ _02521_ VPWR VGND _02522_ sg13g2_buf_1
X_21522_ \atbs_core_0.spike_memory_0.n2398_o[14]\ \atbs_core_0.spike_memory_0.n2397_o[14]\ _02522_ VPWR VGND _01707_ sg13g2_mux2_1
X_21523_ \atbs_core_0.spike_memory_0.n2398_o[15]\ \atbs_core_0.spike_memory_0.n2397_o[15]\ _02522_ VPWR VGND _01708_ sg13g2_mux2_1
X_21524_ \atbs_core_0.spike_memory_0.n2398_o[16]\ \atbs_core_0.spike_memory_0.n2397_o[16]\ _02522_ VPWR VGND _01709_ sg13g2_mux2_1
X_21525_ \atbs_core_0.spike_memory_0.n2398_o[17]\ \atbs_core_0.spike_memory_0.n2397_o[17]\ _02522_ VPWR VGND _01710_ sg13g2_mux2_1
X_21526_ \atbs_core_0.spike_memory_0.n2398_o[18]\ \atbs_core_0.spike_memory_0.n2397_o[18]\ _02522_ VPWR VGND _01711_ sg13g2_mux2_1
X_21527_ \atbs_core_0.spike_memory_0.n2399_o[0]\ VPWR VGND _02523_ sg13g2_buf_1
X_21528_ _02523_ \atbs_core_0.spike_memory_0.n2398_o[0]\ _02522_ VPWR VGND _01712_ sg13g2_mux2_1
X_21529_ \atbs_core_0.spike_memory_0.n2362_o[1]\ \atbs_core_0.spike_memory_0.n2361_o[1]\ _02522_ VPWR VGND _01713_ sg13g2_mux2_1
X_21530_ \atbs_core_0.spike_memory_0.n2399_o[1]\ VPWR VGND _02524_ sg13g2_buf_1
X_21531_ _02524_ \atbs_core_0.spike_memory_0.n2398_o[1]\ _02522_ VPWR VGND _01714_ sg13g2_mux2_1
X_21532_ \atbs_core_0.spike_memory_0.n2399_o[2]\ VPWR VGND _02525_ sg13g2_buf_1
X_21533_ _02525_ \atbs_core_0.spike_memory_0.n2398_o[2]\ _02522_ VPWR VGND _01715_ sg13g2_mux2_1
X_21534_ \atbs_core_0.spike_memory_0.n2399_o[3]\ VPWR VGND _02526_ sg13g2_buf_1
X_21535_ _02526_ \atbs_core_0.spike_memory_0.n2398_o[3]\ _02522_ VPWR VGND _01716_ sg13g2_mux2_1
X_21536_ \atbs_core_0.spike_memory_0.n2399_o[4]\ VPWR VGND _02527_ sg13g2_buf_1
X_21537_ _02521_ VPWR VGND _02528_ sg13g2_buf_1
X_21538_ _02527_ \atbs_core_0.spike_memory_0.n2398_o[4]\ _02528_ VPWR VGND _01717_ sg13g2_mux2_1
X_21539_ \atbs_core_0.spike_memory_0.n2399_o[5]\ VPWR VGND _02529_ sg13g2_buf_1
X_21540_ _02529_ \atbs_core_0.spike_memory_0.n2398_o[5]\ _02528_ VPWR VGND _01718_ sg13g2_mux2_1
X_21541_ \atbs_core_0.spike_memory_0.n2399_o[6]\ VPWR VGND _02530_ sg13g2_buf_1
X_21542_ _02530_ \atbs_core_0.spike_memory_0.n2398_o[6]\ _02528_ VPWR VGND _01719_ sg13g2_mux2_1
X_21543_ \atbs_core_0.spike_memory_0.n2399_o[7]\ VPWR VGND _02531_ sg13g2_buf_1
X_21544_ _02531_ \atbs_core_0.spike_memory_0.n2398_o[7]\ _02528_ VPWR VGND _01720_ sg13g2_mux2_1
X_21545_ \atbs_core_0.spike_memory_0.n2399_o[8]\ VPWR VGND _02532_ sg13g2_buf_1
X_21546_ _02532_ \atbs_core_0.spike_memory_0.n2398_o[8]\ _02528_ VPWR VGND _01721_ sg13g2_mux2_1
X_21547_ \atbs_core_0.spike_memory_0.n2399_o[9]\ VPWR VGND _02533_ sg13g2_buf_1
X_21548_ _02533_ \atbs_core_0.spike_memory_0.n2398_o[9]\ _02528_ VPWR VGND _01722_ sg13g2_mux2_1
X_21549_ \atbs_core_0.spike_memory_0.n2399_o[10]\ VPWR VGND _02534_ sg13g2_buf_1
X_21550_ _02534_ \atbs_core_0.spike_memory_0.n2398_o[10]\ _02528_ VPWR VGND _01723_ sg13g2_mux2_1
X_21551_ \atbs_core_0.spike_memory_0.n2362_o[2]\ \atbs_core_0.spike_memory_0.n2361_o[2]\ _02528_ VPWR VGND _01724_ sg13g2_mux2_1
X_21552_ \atbs_core_0.spike_memory_0.n2399_o[11]\ VPWR VGND _02535_ sg13g2_buf_1
X_21553_ _02535_ \atbs_core_0.spike_memory_0.n2398_o[11]\ _02528_ VPWR VGND _01725_ sg13g2_mux2_1
X_21554_ \atbs_core_0.spike_memory_0.n2399_o[12]\ VPWR VGND _02536_ sg13g2_buf_1
X_21555_ _02536_ \atbs_core_0.spike_memory_0.n2398_o[12]\ _02528_ VPWR VGND _01726_ sg13g2_mux2_1
X_21556_ \atbs_core_0.spike_memory_0.n2399_o[13]\ VPWR VGND _02537_ sg13g2_buf_1
X_21557_ _02521_ VPWR VGND _02538_ sg13g2_buf_1
X_21558_ _02537_ \atbs_core_0.spike_memory_0.n2398_o[13]\ _02538_ VPWR VGND _01727_ sg13g2_mux2_1
X_21559_ \atbs_core_0.spike_memory_0.n2399_o[14]\ VPWR VGND _02539_ sg13g2_buf_1
X_21560_ _02539_ \atbs_core_0.spike_memory_0.n2398_o[14]\ _02538_ VPWR VGND _01728_ sg13g2_mux2_1
X_21561_ \atbs_core_0.spike_memory_0.n2399_o[15]\ VPWR VGND _02540_ sg13g2_buf_1
X_21562_ _02540_ \atbs_core_0.spike_memory_0.n2398_o[15]\ _02538_ VPWR VGND _01729_ sg13g2_mux2_1
X_21563_ \atbs_core_0.spike_memory_0.n2399_o[16]\ VPWR VGND _02541_ sg13g2_buf_1
X_21564_ _02541_ \atbs_core_0.spike_memory_0.n2398_o[16]\ _02538_ VPWR VGND _01730_ sg13g2_mux2_1
X_21565_ \atbs_core_0.spike_memory_0.n2399_o[17]\ VPWR VGND _02542_ sg13g2_buf_1
X_21566_ _02542_ \atbs_core_0.spike_memory_0.n2398_o[17]\ _02538_ VPWR VGND _01731_ sg13g2_mux2_1
X_21567_ \atbs_core_0.spike_memory_0.n2399_o[18]\ VPWR VGND _02543_ sg13g2_buf_1
X_21568_ _02543_ \atbs_core_0.spike_memory_0.n2398_o[18]\ _02538_ VPWR VGND _01732_ sg13g2_mux2_1
X_21569_ \atbs_core_0.spike_memory_0.n2400_o[0]\ VPWR VGND _02544_ sg13g2_buf_1
X_21570_ _02544_ _02523_ _02538_ VPWR VGND _01733_ sg13g2_mux2_1
X_21571_ \atbs_core_0.spike_memory_0.n2400_o[1]\ VPWR VGND _02545_ sg13g2_buf_1
X_21572_ _02545_ _02524_ _02538_ VPWR VGND _01734_ sg13g2_mux2_1
X_21573_ \atbs_core_0.spike_memory_0.n2362_o[3]\ \atbs_core_0.spike_memory_0.n2361_o[3]\ _02538_ VPWR VGND _01735_ sg13g2_mux2_1
X_21574_ \atbs_core_0.spike_memory_0.n2358_o[7]\ \atbs_core_0.spike_memory_0.a_data[7]\ _02538_ VPWR VGND _01736_ sg13g2_mux2_1
X_21575_ \atbs_core_0.spike_memory_0.n2400_o[2]\ VPWR VGND _02546_ sg13g2_buf_1
X_21576_ _02521_ VPWR VGND _02547_ sg13g2_buf_1
X_21577_ _02546_ _02525_ _02547_ VPWR VGND _01737_ sg13g2_mux2_1
X_21578_ \atbs_core_0.spike_memory_0.n2400_o[3]\ VPWR VGND _02548_ sg13g2_buf_1
X_21579_ _02548_ _02526_ _02547_ VPWR VGND _01738_ sg13g2_mux2_1
X_21580_ \atbs_core_0.spike_memory_0.n2400_o[4]\ VPWR VGND _02549_ sg13g2_buf_1
X_21581_ _02549_ _02527_ _02547_ VPWR VGND _01739_ sg13g2_mux2_1
X_21582_ \atbs_core_0.spike_memory_0.n2400_o[5]\ VPWR VGND _02550_ sg13g2_buf_1
X_21583_ _02550_ _02529_ _02547_ VPWR VGND _01740_ sg13g2_mux2_1
X_21584_ \atbs_core_0.spike_memory_0.n2400_o[6]\ VPWR VGND _02551_ sg13g2_buf_1
X_21585_ _02551_ _02530_ _02547_ VPWR VGND _01741_ sg13g2_mux2_1
X_21586_ \atbs_core_0.spike_memory_0.n2400_o[7]\ VPWR VGND _02552_ sg13g2_buf_1
X_21587_ _02552_ _02531_ _02547_ VPWR VGND _01742_ sg13g2_mux2_1
X_21588_ \atbs_core_0.spike_memory_0.n2400_o[8]\ VPWR VGND _02553_ sg13g2_buf_1
X_21589_ _02553_ _02532_ _02547_ VPWR VGND _01743_ sg13g2_mux2_1
X_21590_ \atbs_core_0.spike_memory_0.n2400_o[9]\ VPWR VGND _02554_ sg13g2_buf_1
X_21591_ _02554_ _02533_ _02547_ VPWR VGND _01744_ sg13g2_mux2_1
X_21592_ \atbs_core_0.spike_memory_0.n2400_o[10]\ VPWR VGND _02555_ sg13g2_buf_1
X_21593_ _02555_ _02534_ _02547_ VPWR VGND _01745_ sg13g2_mux2_1
X_21594_ \atbs_core_0.spike_memory_0.n2400_o[11]\ VPWR VGND _02556_ sg13g2_buf_1
X_21595_ _02556_ _02535_ _02547_ VPWR VGND _01746_ sg13g2_mux2_1
X_21596_ _02521_ VPWR VGND _02557_ sg13g2_buf_1
X_21597_ \atbs_core_0.spike_memory_0.n2362_o[4]\ \atbs_core_0.spike_memory_0.n2361_o[4]\ _02557_ VPWR VGND _01747_ sg13g2_mux2_1
X_21598_ \atbs_core_0.spike_memory_0.n2400_o[12]\ VPWR VGND _02558_ sg13g2_buf_1
X_21599_ _02558_ _02536_ _02557_ VPWR VGND _01748_ sg13g2_mux2_1
X_21600_ \atbs_core_0.spike_memory_0.n2400_o[13]\ VPWR VGND _02559_ sg13g2_buf_1
X_21601_ _02559_ _02537_ _02557_ VPWR VGND _01749_ sg13g2_mux2_1
X_21602_ \atbs_core_0.spike_memory_0.n2400_o[14]\ VPWR VGND _02560_ sg13g2_buf_1
X_21603_ _02560_ _02539_ _02557_ VPWR VGND _01750_ sg13g2_mux2_1
X_21604_ \atbs_core_0.spike_memory_0.n2400_o[15]\ VPWR VGND _02561_ sg13g2_buf_1
X_21605_ _02561_ _02540_ _02557_ VPWR VGND _01751_ sg13g2_mux2_1
X_21606_ \atbs_core_0.spike_memory_0.n2400_o[16]\ VPWR VGND _02562_ sg13g2_buf_1
X_21607_ _02562_ _02541_ _02557_ VPWR VGND _01752_ sg13g2_mux2_1
X_21608_ \atbs_core_0.spike_memory_0.n2400_o[17]\ VPWR VGND _02563_ sg13g2_buf_1
X_21609_ _02563_ _02542_ _02557_ VPWR VGND _01753_ sg13g2_mux2_1
X_21610_ \atbs_core_0.spike_memory_0.n2400_o[18]\ VPWR VGND _02564_ sg13g2_buf_1
X_21611_ _02564_ _02543_ _02557_ VPWR VGND _01754_ sg13g2_mux2_1
X_21612_ \atbs_core_0.spike_memory_0.n2401_o[0]\ _02544_ _02557_ VPWR VGND _01755_ sg13g2_mux2_1
X_21613_ \atbs_core_0.spike_memory_0.n2401_o[1]\ _02545_ _02557_ VPWR VGND _01756_ sg13g2_mux2_1
X_21614_ _02521_ VPWR VGND _02565_ sg13g2_buf_1
X_21615_ \atbs_core_0.spike_memory_0.n2401_o[2]\ _02546_ _02565_ VPWR VGND _01757_ sg13g2_mux2_1
X_21616_ \atbs_core_0.spike_memory_0.n2362_o[5]\ \atbs_core_0.spike_memory_0.n2361_o[5]\ _02565_ VPWR VGND _01758_ sg13g2_mux2_1
X_21617_ \atbs_core_0.spike_memory_0.n2401_o[3]\ _02548_ _02565_ VPWR VGND _01759_ sg13g2_mux2_1
X_21618_ \atbs_core_0.spike_memory_0.n2401_o[4]\ _02549_ _02565_ VPWR VGND _01760_ sg13g2_mux2_1
X_21619_ \atbs_core_0.spike_memory_0.n2401_o[5]\ _02550_ _02565_ VPWR VGND _01761_ sg13g2_mux2_1
X_21620_ \atbs_core_0.spike_memory_0.n2401_o[6]\ _02551_ _02565_ VPWR VGND _01762_ sg13g2_mux2_1
X_21621_ \atbs_core_0.spike_memory_0.n2401_o[7]\ _02552_ _02565_ VPWR VGND _01763_ sg13g2_mux2_1
X_21622_ \atbs_core_0.spike_memory_0.n2401_o[8]\ _02553_ _02565_ VPWR VGND _01764_ sg13g2_mux2_1
X_21623_ \atbs_core_0.spike_memory_0.n2401_o[9]\ _02554_ _02565_ VPWR VGND _01765_ sg13g2_mux2_1
X_21624_ \atbs_core_0.spike_memory_0.n2401_o[10]\ _02555_ _02565_ VPWR VGND _01766_ sg13g2_mux2_1
X_21625_ _02521_ VPWR VGND _02566_ sg13g2_buf_1
X_21626_ \atbs_core_0.spike_memory_0.n2401_o[11]\ _02556_ _02566_ VPWR VGND _01767_ sg13g2_mux2_1
X_21627_ \atbs_core_0.spike_memory_0.n2401_o[12]\ _02558_ _02566_ VPWR VGND _01768_ sg13g2_mux2_1
X_21628_ \atbs_core_0.spike_memory_0.n2362_o[6]\ \atbs_core_0.spike_memory_0.n2361_o[6]\ _02566_ VPWR VGND _01769_ sg13g2_mux2_1
X_21629_ \atbs_core_0.spike_memory_0.n2401_o[13]\ _02559_ _02566_ VPWR VGND _01770_ sg13g2_mux2_1
X_21630_ \atbs_core_0.spike_memory_0.n2401_o[14]\ _02560_ _02566_ VPWR VGND _01771_ sg13g2_mux2_1
X_21631_ \atbs_core_0.spike_memory_0.n2401_o[15]\ _02561_ _02566_ VPWR VGND _01772_ sg13g2_mux2_1
X_21632_ \atbs_core_0.spike_memory_0.n2401_o[16]\ _02562_ _02566_ VPWR VGND _01773_ sg13g2_mux2_1
X_21633_ \atbs_core_0.spike_memory_0.n2401_o[17]\ _02563_ _02566_ VPWR VGND _01774_ sg13g2_mux2_1
X_21634_ \atbs_core_0.spike_memory_0.n2401_o[18]\ _02564_ _02566_ VPWR VGND _01775_ sg13g2_mux2_1
X_21635_ \atbs_core_0.spike_memory_0.n2402_o[0]\ \atbs_core_0.spike_memory_0.n2401_o[0]\ _02566_ VPWR VGND _01776_ sg13g2_mux2_1
X_21636_ _12511_ VPWR VGND _02567_ sg13g2_buf_1
X_21637_ _02567_ VPWR VGND _02568_ sg13g2_buf_1
X_21638_ \atbs_core_0.spike_memory_0.n2402_o[1]\ \atbs_core_0.spike_memory_0.n2401_o[1]\ _02568_ VPWR VGND _01777_ sg13g2_mux2_1
X_21639_ \atbs_core_0.spike_memory_0.n2402_o[2]\ \atbs_core_0.spike_memory_0.n2401_o[2]\ _02568_ VPWR VGND _01778_ sg13g2_mux2_1
X_21640_ \atbs_core_0.spike_memory_0.n2402_o[3]\ \atbs_core_0.spike_memory_0.n2401_o[3]\ _02568_ VPWR VGND _01779_ sg13g2_mux2_1
X_21641_ \atbs_core_0.spike_memory_0.n2362_o[7]\ \atbs_core_0.spike_memory_0.n2361_o[7]\ _02568_ VPWR VGND _01780_ sg13g2_mux2_1
X_21642_ \atbs_core_0.spike_memory_0.n2402_o[4]\ \atbs_core_0.spike_memory_0.n2401_o[4]\ _02568_ VPWR VGND _01781_ sg13g2_mux2_1
X_21643_ \atbs_core_0.spike_memory_0.n2402_o[5]\ \atbs_core_0.spike_memory_0.n2401_o[5]\ _02568_ VPWR VGND _01782_ sg13g2_mux2_1
X_21644_ \atbs_core_0.spike_memory_0.n2402_o[6]\ \atbs_core_0.spike_memory_0.n2401_o[6]\ _02568_ VPWR VGND _01783_ sg13g2_mux2_1
X_21645_ \atbs_core_0.spike_memory_0.n2402_o[7]\ \atbs_core_0.spike_memory_0.n2401_o[7]\ _02568_ VPWR VGND _01784_ sg13g2_mux2_1
X_21646_ \atbs_core_0.spike_memory_0.n2402_o[8]\ \atbs_core_0.spike_memory_0.n2401_o[8]\ _02568_ VPWR VGND _01785_ sg13g2_mux2_1
X_21647_ \atbs_core_0.spike_memory_0.n2402_o[9]\ \atbs_core_0.spike_memory_0.n2401_o[9]\ _02568_ VPWR VGND _01786_ sg13g2_mux2_1
X_21648_ _02567_ VPWR VGND _02569_ sg13g2_buf_1
X_21649_ \atbs_core_0.spike_memory_0.n2402_o[10]\ \atbs_core_0.spike_memory_0.n2401_o[10]\ _02569_ VPWR VGND _01787_ sg13g2_mux2_1
X_21650_ \atbs_core_0.spike_memory_0.n2402_o[11]\ \atbs_core_0.spike_memory_0.n2401_o[11]\ _02569_ VPWR VGND _01788_ sg13g2_mux2_1
X_21651_ \atbs_core_0.spike_memory_0.n2402_o[12]\ \atbs_core_0.spike_memory_0.n2401_o[12]\ _02569_ VPWR VGND _01789_ sg13g2_mux2_1
X_21652_ \atbs_core_0.spike_memory_0.n2402_o[13]\ \atbs_core_0.spike_memory_0.n2401_o[13]\ _02569_ VPWR VGND _01790_ sg13g2_mux2_1
X_21653_ \atbs_core_0.spike_memory_0.n2362_o[8]\ \atbs_core_0.spike_memory_0.n2361_o[8]\ _02569_ VPWR VGND _01791_ sg13g2_mux2_1
X_21654_ \atbs_core_0.spike_memory_0.n2402_o[14]\ \atbs_core_0.spike_memory_0.n2401_o[14]\ _02569_ VPWR VGND _01792_ sg13g2_mux2_1
X_21655_ \atbs_core_0.spike_memory_0.n2402_o[15]\ \atbs_core_0.spike_memory_0.n2401_o[15]\ _02569_ VPWR VGND _01793_ sg13g2_mux2_1
X_21656_ \atbs_core_0.spike_memory_0.n2402_o[16]\ \atbs_core_0.spike_memory_0.n2401_o[16]\ _02569_ VPWR VGND _01794_ sg13g2_mux2_1
X_21657_ \atbs_core_0.spike_memory_0.n2402_o[17]\ \atbs_core_0.spike_memory_0.n2401_o[17]\ _02569_ VPWR VGND _01795_ sg13g2_mux2_1
X_21658_ \atbs_core_0.spike_memory_0.n2402_o[18]\ \atbs_core_0.spike_memory_0.n2401_o[18]\ _02569_ VPWR VGND _01796_ sg13g2_mux2_1
X_21659_ \atbs_core_0.spike_memory_0.n2403_o[0]\ VPWR VGND _02570_ sg13g2_buf_1
X_21660_ _02567_ VPWR VGND _02571_ sg13g2_buf_1
X_21661_ _02570_ \atbs_core_0.spike_memory_0.n2402_o[0]\ _02571_ VPWR VGND _01797_ sg13g2_mux2_1
X_21662_ \atbs_core_0.spike_memory_0.n2403_o[1]\ VPWR VGND _02572_ sg13g2_buf_1
X_21663_ _02572_ \atbs_core_0.spike_memory_0.n2402_o[1]\ _02571_ VPWR VGND _01798_ sg13g2_mux2_1
X_21664_ \atbs_core_0.spike_memory_0.n2403_o[2]\ VPWR VGND _02573_ sg13g2_buf_1
X_21665_ _02573_ \atbs_core_0.spike_memory_0.n2402_o[2]\ _02571_ VPWR VGND _01799_ sg13g2_mux2_1
X_21666_ \atbs_core_0.spike_memory_0.n2403_o[3]\ VPWR VGND _02574_ sg13g2_buf_1
X_21667_ _02574_ \atbs_core_0.spike_memory_0.n2402_o[3]\ _02571_ VPWR VGND _01800_ sg13g2_mux2_1
X_21668_ \atbs_core_0.spike_memory_0.n2403_o[4]\ VPWR VGND _02575_ sg13g2_buf_1
X_21669_ _02575_ \atbs_core_0.spike_memory_0.n2402_o[4]\ _02571_ VPWR VGND _01801_ sg13g2_mux2_1
X_21670_ \atbs_core_0.spike_memory_0.n2362_o[9]\ \atbs_core_0.spike_memory_0.n2361_o[9]\ _02571_ VPWR VGND _01802_ sg13g2_mux2_1
X_21671_ \atbs_core_0.spike_memory_0.n2403_o[5]\ VPWR VGND _02576_ sg13g2_buf_1
X_21672_ _02576_ \atbs_core_0.spike_memory_0.n2402_o[5]\ _02571_ VPWR VGND _01803_ sg13g2_mux2_1
X_21673_ \atbs_core_0.spike_memory_0.n2403_o[6]\ VPWR VGND _02577_ sg13g2_buf_1
X_21674_ _02577_ \atbs_core_0.spike_memory_0.n2402_o[6]\ _02571_ VPWR VGND _01804_ sg13g2_mux2_1
X_21675_ \atbs_core_0.spike_memory_0.n2403_o[7]\ VPWR VGND _02578_ sg13g2_buf_1
X_21676_ _02578_ \atbs_core_0.spike_memory_0.n2402_o[7]\ _02571_ VPWR VGND _01805_ sg13g2_mux2_1
X_21677_ \atbs_core_0.spike_memory_0.n2403_o[8]\ VPWR VGND _02579_ sg13g2_buf_1
X_21678_ _02579_ \atbs_core_0.spike_memory_0.n2402_o[8]\ _02571_ VPWR VGND _01806_ sg13g2_mux2_1
X_21679_ \atbs_core_0.spike_memory_0.n2403_o[9]\ VPWR VGND _02580_ sg13g2_buf_1
X_21680_ _02567_ VPWR VGND _02581_ sg13g2_buf_1
X_21681_ _02580_ \atbs_core_0.spike_memory_0.n2402_o[9]\ _02581_ VPWR VGND _01807_ sg13g2_mux2_1
X_21682_ \atbs_core_0.spike_memory_0.n2403_o[10]\ VPWR VGND _02582_ sg13g2_buf_1
X_21683_ _02582_ \atbs_core_0.spike_memory_0.n2402_o[10]\ _02581_ VPWR VGND _01808_ sg13g2_mux2_1
X_21684_ \atbs_core_0.spike_memory_0.n2403_o[11]\ VPWR VGND _02583_ sg13g2_buf_1
X_21685_ _02583_ \atbs_core_0.spike_memory_0.n2402_o[11]\ _02581_ VPWR VGND _01809_ sg13g2_mux2_1
X_21686_ \atbs_core_0.spike_memory_0.n2403_o[12]\ VPWR VGND _02584_ sg13g2_buf_1
X_21687_ _02584_ \atbs_core_0.spike_memory_0.n2402_o[12]\ _02581_ VPWR VGND _01810_ sg13g2_mux2_1
X_21688_ \atbs_core_0.spike_memory_0.n2403_o[13]\ VPWR VGND _02585_ sg13g2_buf_1
X_21689_ _02585_ \atbs_core_0.spike_memory_0.n2402_o[13]\ _02581_ VPWR VGND _01811_ sg13g2_mux2_1
X_21690_ \atbs_core_0.spike_memory_0.n2403_o[14]\ VPWR VGND _02586_ sg13g2_buf_1
X_21691_ _02586_ \atbs_core_0.spike_memory_0.n2402_o[14]\ _02581_ VPWR VGND _01812_ sg13g2_mux2_1
X_21692_ \atbs_core_0.spike_memory_0.n2362_o[10]\ \atbs_core_0.spike_memory_0.n2361_o[10]\ _02581_ VPWR VGND _01813_ sg13g2_mux2_1
X_21693_ \atbs_core_0.spike_memory_0.n2403_o[15]\ VPWR VGND _02587_ sg13g2_buf_1
X_21694_ _02587_ \atbs_core_0.spike_memory_0.n2402_o[15]\ _02581_ VPWR VGND _01814_ sg13g2_mux2_1
X_21695_ \atbs_core_0.spike_memory_0.n2403_o[16]\ VPWR VGND _02588_ sg13g2_buf_1
X_21696_ _02588_ \atbs_core_0.spike_memory_0.n2402_o[16]\ _02581_ VPWR VGND _01815_ sg13g2_mux2_1
X_21697_ \atbs_core_0.spike_memory_0.n2403_o[17]\ VPWR VGND _02589_ sg13g2_buf_1
X_21698_ _02589_ \atbs_core_0.spike_memory_0.n2402_o[17]\ _02581_ VPWR VGND _01816_ sg13g2_mux2_1
X_21699_ \atbs_core_0.spike_memory_0.n2403_o[18]\ VPWR VGND _02590_ sg13g2_buf_1
X_21700_ _02567_ VPWR VGND _02591_ sg13g2_buf_1
X_21701_ _02590_ \atbs_core_0.spike_memory_0.n2402_o[18]\ _02591_ VPWR VGND _01817_ sg13g2_mux2_1
X_21702_ \atbs_core_0.spike_memory_0.n2404_o[0]\ VPWR VGND _02592_ sg13g2_buf_1
X_21703_ _02592_ _02570_ _02591_ VPWR VGND _01818_ sg13g2_mux2_1
X_21704_ \atbs_core_0.spike_memory_0.n2404_o[1]\ VPWR VGND _02593_ sg13g2_buf_1
X_21705_ _02593_ _02572_ _02591_ VPWR VGND _01819_ sg13g2_mux2_1
X_21706_ \atbs_core_0.spike_memory_0.n2404_o[2]\ VPWR VGND _02594_ sg13g2_buf_1
X_21707_ _02594_ _02573_ _02591_ VPWR VGND _01820_ sg13g2_mux2_1
X_21708_ \atbs_core_0.spike_memory_0.n2404_o[3]\ VPWR VGND _02595_ sg13g2_buf_1
X_21709_ _02595_ _02574_ _02591_ VPWR VGND _01821_ sg13g2_mux2_1
X_21710_ \atbs_core_0.spike_memory_0.n2404_o[4]\ VPWR VGND _02596_ sg13g2_buf_1
X_21711_ _02596_ _02575_ _02591_ VPWR VGND _01822_ sg13g2_mux2_1
X_21712_ \atbs_core_0.spike_memory_0.n2404_o[5]\ VPWR VGND _02597_ sg13g2_buf_1
X_21713_ _02597_ _02576_ _02591_ VPWR VGND _01823_ sg13g2_mux2_1
X_21714_ \atbs_core_0.spike_memory_0.n2362_o[11]\ \atbs_core_0.spike_memory_0.n2361_o[11]\ _02591_ VPWR VGND _01824_ sg13g2_mux2_1
X_21715_ \atbs_core_0.spike_memory_0.n2404_o[6]\ VPWR VGND _02598_ sg13g2_buf_1
X_21716_ _02598_ _02577_ _02591_ VPWR VGND _01825_ sg13g2_mux2_1
X_21717_ \atbs_core_0.spike_memory_0.n2404_o[7]\ VPWR VGND _02599_ sg13g2_buf_1
X_21718_ _02599_ _02578_ _02591_ VPWR VGND _01826_ sg13g2_mux2_1
X_21719_ \atbs_core_0.spike_memory_0.n2404_o[8]\ VPWR VGND _02600_ sg13g2_buf_1
X_21720_ _02567_ VPWR VGND _02601_ sg13g2_buf_1
X_21721_ _02600_ _02579_ _02601_ VPWR VGND _01827_ sg13g2_mux2_1
X_21722_ \atbs_core_0.spike_memory_0.n2404_o[9]\ VPWR VGND _02602_ sg13g2_buf_1
X_21723_ _02602_ _02580_ _02601_ VPWR VGND _01828_ sg13g2_mux2_1
X_21724_ \atbs_core_0.spike_memory_0.n2404_o[10]\ VPWR VGND _02603_ sg13g2_buf_1
X_21725_ _02603_ _02582_ _02601_ VPWR VGND _01829_ sg13g2_mux2_1
X_21726_ \atbs_core_0.spike_memory_0.n2404_o[11]\ VPWR VGND _02604_ sg13g2_buf_1
X_21727_ _02604_ _02583_ _02601_ VPWR VGND _01830_ sg13g2_mux2_1
X_21728_ \atbs_core_0.spike_memory_0.n2404_o[12]\ VPWR VGND _02605_ sg13g2_buf_1
X_21729_ _02605_ _02584_ _02601_ VPWR VGND _01831_ sg13g2_mux2_1
X_21730_ \atbs_core_0.spike_memory_0.n2404_o[13]\ VPWR VGND _02606_ sg13g2_buf_1
X_21731_ _02606_ _02585_ _02601_ VPWR VGND _01832_ sg13g2_mux2_1
X_21732_ \atbs_core_0.spike_memory_0.n2404_o[14]\ VPWR VGND _02607_ sg13g2_buf_1
X_21733_ _02607_ _02586_ _02601_ VPWR VGND _01833_ sg13g2_mux2_1
X_21734_ \atbs_core_0.spike_memory_0.n2404_o[15]\ VPWR VGND _02608_ sg13g2_buf_1
X_21735_ _02608_ _02587_ _02601_ VPWR VGND _01834_ sg13g2_mux2_1
X_21736_ \atbs_core_0.spike_memory_0.n2362_o[12]\ \atbs_core_0.spike_memory_0.n2361_o[12]\ _02601_ VPWR VGND _01835_ sg13g2_mux2_1
X_21737_ \atbs_core_0.spike_memory_0.n2404_o[16]\ VPWR VGND _02609_ sg13g2_buf_1
X_21738_ _02609_ _02588_ _02601_ VPWR VGND _01836_ sg13g2_mux2_1
X_21739_ \atbs_core_0.spike_memory_0.n2404_o[17]\ VPWR VGND _02610_ sg13g2_buf_1
X_21740_ _02567_ VPWR VGND _02611_ sg13g2_buf_1
X_21741_ _02610_ _02589_ _02611_ VPWR VGND _01837_ sg13g2_mux2_1
X_21742_ \atbs_core_0.spike_memory_0.n2404_o[18]\ VPWR VGND _02612_ sg13g2_buf_1
X_21743_ _02612_ _02590_ _02611_ VPWR VGND _01838_ sg13g2_mux2_1
X_21744_ \atbs_core_0.spike_memory_0.n2405_o[0]\ _02592_ _02611_ VPWR VGND _01839_ sg13g2_mux2_1
X_21745_ \atbs_core_0.spike_memory_0.n2405_o[1]\ _02593_ _02611_ VPWR VGND _01840_ sg13g2_mux2_1
X_21746_ \atbs_core_0.spike_memory_0.n2405_o[2]\ _02594_ _02611_ VPWR VGND _01841_ sg13g2_mux2_1
X_21747_ \atbs_core_0.spike_memory_0.n2405_o[3]\ _02595_ _02611_ VPWR VGND _01842_ sg13g2_mux2_1
X_21748_ \atbs_core_0.spike_memory_0.n2405_o[4]\ _02596_ _02611_ VPWR VGND _01843_ sg13g2_mux2_1
X_21749_ \atbs_core_0.spike_memory_0.n2405_o[5]\ _02597_ _02611_ VPWR VGND _01844_ sg13g2_mux2_1
X_21750_ \atbs_core_0.spike_memory_0.n2405_o[6]\ _02598_ _02611_ VPWR VGND _01845_ sg13g2_mux2_1
X_21751_ \atbs_core_0.spike_memory_0.n2362_o[13]\ \atbs_core_0.spike_memory_0.n2361_o[13]\ _02611_ VPWR VGND _01846_ sg13g2_mux2_1
X_21752_ _12511_ VPWR VGND _02613_ sg13g2_buf_1
X_21753_ _02613_ VPWR VGND _02614_ sg13g2_buf_1
X_21754_ \atbs_core_0.spike_memory_0.n2358_o[8]\ \atbs_core_0.spike_memory_0.a_data[8]\ _02614_ VPWR VGND _01847_ sg13g2_mux2_1
X_21755_ \atbs_core_0.spike_memory_0.n2405_o[7]\ _02599_ _02614_ VPWR VGND _01848_ sg13g2_mux2_1
X_21756_ \atbs_core_0.spike_memory_0.n2405_o[8]\ _02600_ _02614_ VPWR VGND _01849_ sg13g2_mux2_1
X_21757_ \atbs_core_0.spike_memory_0.n2405_o[9]\ _02602_ _02614_ VPWR VGND _01850_ sg13g2_mux2_1
X_21758_ \atbs_core_0.spike_memory_0.n2405_o[10]\ _02603_ _02614_ VPWR VGND _01851_ sg13g2_mux2_1
X_21759_ \atbs_core_0.spike_memory_0.n2405_o[11]\ _02604_ _02614_ VPWR VGND _01852_ sg13g2_mux2_1
X_21760_ \atbs_core_0.spike_memory_0.n2405_o[12]\ _02605_ _02614_ VPWR VGND _01853_ sg13g2_mux2_1
X_21761_ \atbs_core_0.spike_memory_0.n2405_o[13]\ _02606_ _02614_ VPWR VGND _01854_ sg13g2_mux2_1
X_21762_ \atbs_core_0.spike_memory_0.n2405_o[14]\ _02607_ _02614_ VPWR VGND _01855_ sg13g2_mux2_1
X_21763_ \atbs_core_0.spike_memory_0.n2405_o[15]\ _02608_ _02614_ VPWR VGND _01856_ sg13g2_mux2_1
X_21764_ _02613_ VPWR VGND _02615_ sg13g2_buf_1
X_21765_ \atbs_core_0.spike_memory_0.n2405_o[16]\ _02609_ _02615_ VPWR VGND _01857_ sg13g2_mux2_1
X_21766_ \atbs_core_0.spike_memory_0.n2362_o[14]\ \atbs_core_0.spike_memory_0.n2361_o[14]\ _02615_ VPWR VGND _01858_ sg13g2_mux2_1
X_21767_ \atbs_core_0.spike_memory_0.n2405_o[17]\ _02610_ _02615_ VPWR VGND _01859_ sg13g2_mux2_1
X_21768_ \atbs_core_0.spike_memory_0.n2405_o[18]\ _02612_ _02615_ VPWR VGND _01860_ sg13g2_mux2_1
X_21769_ \atbs_core_0.spike_memory_0.n2406_o[0]\ \atbs_core_0.spike_memory_0.n2405_o[0]\ _02615_ VPWR VGND _01861_ sg13g2_mux2_1
X_21770_ \atbs_core_0.spike_memory_0.n2406_o[1]\ \atbs_core_0.spike_memory_0.n2405_o[1]\ _02615_ VPWR VGND _01862_ sg13g2_mux2_1
X_21771_ \atbs_core_0.spike_memory_0.n2406_o[2]\ \atbs_core_0.spike_memory_0.n2405_o[2]\ _02615_ VPWR VGND _01863_ sg13g2_mux2_1
X_21772_ \atbs_core_0.spike_memory_0.n2406_o[3]\ \atbs_core_0.spike_memory_0.n2405_o[3]\ _02615_ VPWR VGND _01864_ sg13g2_mux2_1
X_21773_ \atbs_core_0.spike_memory_0.n2406_o[4]\ \atbs_core_0.spike_memory_0.n2405_o[4]\ _02615_ VPWR VGND _01865_ sg13g2_mux2_1
X_21774_ \atbs_core_0.spike_memory_0.n2406_o[5]\ \atbs_core_0.spike_memory_0.n2405_o[5]\ _02615_ VPWR VGND _01866_ sg13g2_mux2_1
X_21775_ _02613_ VPWR VGND _02616_ sg13g2_buf_1
X_21776_ \atbs_core_0.spike_memory_0.n2406_o[6]\ \atbs_core_0.spike_memory_0.n2405_o[6]\ _02616_ VPWR VGND _01867_ sg13g2_mux2_1
X_21777_ \atbs_core_0.spike_memory_0.n2406_o[7]\ \atbs_core_0.spike_memory_0.n2405_o[7]\ _02616_ VPWR VGND _01868_ sg13g2_mux2_1
X_21778_ \atbs_core_0.spike_memory_0.n2362_o[15]\ \atbs_core_0.spike_memory_0.n2361_o[15]\ _02616_ VPWR VGND _01869_ sg13g2_mux2_1
X_21779_ \atbs_core_0.spike_memory_0.n2406_o[8]\ \atbs_core_0.spike_memory_0.n2405_o[8]\ _02616_ VPWR VGND _01870_ sg13g2_mux2_1
X_21780_ \atbs_core_0.spike_memory_0.n2406_o[9]\ \atbs_core_0.spike_memory_0.n2405_o[9]\ _02616_ VPWR VGND _01871_ sg13g2_mux2_1
X_21781_ \atbs_core_0.spike_memory_0.n2406_o[10]\ \atbs_core_0.spike_memory_0.n2405_o[10]\ _02616_ VPWR VGND _01872_ sg13g2_mux2_1
X_21782_ \atbs_core_0.spike_memory_0.n2406_o[11]\ \atbs_core_0.spike_memory_0.n2405_o[11]\ _02616_ VPWR VGND _01873_ sg13g2_mux2_1
X_21783_ \atbs_core_0.spike_memory_0.n2406_o[12]\ \atbs_core_0.spike_memory_0.n2405_o[12]\ _02616_ VPWR VGND _01874_ sg13g2_mux2_1
X_21784_ \atbs_core_0.spike_memory_0.n2406_o[13]\ \atbs_core_0.spike_memory_0.n2405_o[13]\ _02616_ VPWR VGND _01875_ sg13g2_mux2_1
X_21785_ \atbs_core_0.spike_memory_0.n2406_o[14]\ \atbs_core_0.spike_memory_0.n2405_o[14]\ _02616_ VPWR VGND _01876_ sg13g2_mux2_1
X_21786_ _02613_ VPWR VGND _02617_ sg13g2_buf_1
X_21787_ \atbs_core_0.spike_memory_0.n2406_o[15]\ \atbs_core_0.spike_memory_0.n2405_o[15]\ _02617_ VPWR VGND _01877_ sg13g2_mux2_1
X_21788_ \atbs_core_0.spike_memory_0.n2406_o[16]\ \atbs_core_0.spike_memory_0.n2405_o[16]\ _02617_ VPWR VGND _01878_ sg13g2_mux2_1
X_21789_ \atbs_core_0.spike_memory_0.n2406_o[17]\ \atbs_core_0.spike_memory_0.n2405_o[17]\ _02617_ VPWR VGND _01879_ sg13g2_mux2_1
X_21790_ \atbs_core_0.spike_memory_0.n2362_o[16]\ \atbs_core_0.spike_memory_0.n2361_o[16]\ _02617_ VPWR VGND _01880_ sg13g2_mux2_1
X_21791_ \atbs_core_0.spike_memory_0.n2406_o[18]\ \atbs_core_0.spike_memory_0.n2405_o[18]\ _02617_ VPWR VGND _01881_ sg13g2_mux2_1
X_21792_ \atbs_core_0.spike_memory_0.n2407_o[0]\ VPWR VGND _02618_ sg13g2_buf_1
X_21793_ _02618_ \atbs_core_0.spike_memory_0.n2406_o[0]\ _02617_ VPWR VGND _01882_ sg13g2_mux2_1
X_21794_ \atbs_core_0.spike_memory_0.n2407_o[1]\ VPWR VGND _02619_ sg13g2_buf_1
X_21795_ _02619_ \atbs_core_0.spike_memory_0.n2406_o[1]\ _02617_ VPWR VGND _01883_ sg13g2_mux2_1
X_21796_ \atbs_core_0.spike_memory_0.n2407_o[2]\ VPWR VGND _02620_ sg13g2_buf_1
X_21797_ _02620_ \atbs_core_0.spike_memory_0.n2406_o[2]\ _02617_ VPWR VGND _01884_ sg13g2_mux2_1
X_21798_ \atbs_core_0.spike_memory_0.n2407_o[3]\ VPWR VGND _02621_ sg13g2_buf_1
X_21799_ _02621_ \atbs_core_0.spike_memory_0.n2406_o[3]\ _02617_ VPWR VGND _01885_ sg13g2_mux2_1
X_21800_ \atbs_core_0.spike_memory_0.n2407_o[4]\ VPWR VGND _02622_ sg13g2_buf_1
X_21801_ _02622_ \atbs_core_0.spike_memory_0.n2406_o[4]\ _02617_ VPWR VGND _01886_ sg13g2_mux2_1
X_21802_ \atbs_core_0.spike_memory_0.n2407_o[5]\ VPWR VGND _02623_ sg13g2_buf_1
X_21803_ _02613_ VPWR VGND _02624_ sg13g2_buf_1
X_21804_ _02623_ \atbs_core_0.spike_memory_0.n2406_o[5]\ _02624_ VPWR VGND _01887_ sg13g2_mux2_1
X_21805_ \atbs_core_0.spike_memory_0.n2407_o[6]\ VPWR VGND _02625_ sg13g2_buf_1
X_21806_ _02625_ \atbs_core_0.spike_memory_0.n2406_o[6]\ _02624_ VPWR VGND _01888_ sg13g2_mux2_1
X_21807_ \atbs_core_0.spike_memory_0.n2407_o[7]\ VPWR VGND _02626_ sg13g2_buf_1
X_21808_ _02626_ \atbs_core_0.spike_memory_0.n2406_o[7]\ _02624_ VPWR VGND _01889_ sg13g2_mux2_1
X_21809_ \atbs_core_0.spike_memory_0.n2407_o[8]\ VPWR VGND _02627_ sg13g2_buf_1
X_21810_ _02627_ \atbs_core_0.spike_memory_0.n2406_o[8]\ _02624_ VPWR VGND _01890_ sg13g2_mux2_1
X_21811_ \atbs_core_0.spike_memory_0.n2362_o[17]\ \atbs_core_0.spike_memory_0.n2361_o[17]\ _02624_ VPWR VGND _01891_ sg13g2_mux2_1
X_21812_ \atbs_core_0.spike_memory_0.n2407_o[9]\ VPWR VGND _02628_ sg13g2_buf_1
X_21813_ _02628_ \atbs_core_0.spike_memory_0.n2406_o[9]\ _02624_ VPWR VGND _01892_ sg13g2_mux2_1
X_21814_ \atbs_core_0.spike_memory_0.n2407_o[10]\ VPWR VGND _02629_ sg13g2_buf_1
X_21815_ _02629_ \atbs_core_0.spike_memory_0.n2406_o[10]\ _02624_ VPWR VGND _01893_ sg13g2_mux2_1
X_21816_ \atbs_core_0.spike_memory_0.n2407_o[11]\ VPWR VGND _02630_ sg13g2_buf_1
X_21817_ _02630_ \atbs_core_0.spike_memory_0.n2406_o[11]\ _02624_ VPWR VGND _01894_ sg13g2_mux2_1
X_21818_ \atbs_core_0.spike_memory_0.n2407_o[12]\ VPWR VGND _02631_ sg13g2_buf_1
X_21819_ _02631_ \atbs_core_0.spike_memory_0.n2406_o[12]\ _02624_ VPWR VGND _01895_ sg13g2_mux2_1
X_21820_ \atbs_core_0.spike_memory_0.n2407_o[13]\ VPWR VGND _02632_ sg13g2_buf_1
X_21821_ _02632_ \atbs_core_0.spike_memory_0.n2406_o[13]\ _02624_ VPWR VGND _01896_ sg13g2_mux2_1
X_21822_ \atbs_core_0.spike_memory_0.n2407_o[14]\ VPWR VGND _02633_ sg13g2_buf_1
X_21823_ _02613_ VPWR VGND _02634_ sg13g2_buf_1
X_21824_ _02633_ \atbs_core_0.spike_memory_0.n2406_o[14]\ _02634_ VPWR VGND _01897_ sg13g2_mux2_1
X_21825_ \atbs_core_0.spike_memory_0.n2407_o[15]\ VPWR VGND _02635_ sg13g2_buf_1
X_21826_ _02635_ \atbs_core_0.spike_memory_0.n2406_o[15]\ _02634_ VPWR VGND _01898_ sg13g2_mux2_1
X_21827_ \atbs_core_0.spike_memory_0.n2407_o[16]\ VPWR VGND _02636_ sg13g2_buf_1
X_21828_ _02636_ \atbs_core_0.spike_memory_0.n2406_o[16]\ _02634_ VPWR VGND _01899_ sg13g2_mux2_1
X_21829_ \atbs_core_0.spike_memory_0.n2407_o[17]\ VPWR VGND _02637_ sg13g2_buf_1
X_21830_ _02637_ \atbs_core_0.spike_memory_0.n2406_o[17]\ _02634_ VPWR VGND _01900_ sg13g2_mux2_1
X_21831_ \atbs_core_0.spike_memory_0.n2407_o[18]\ VPWR VGND _02638_ sg13g2_buf_1
X_21832_ _02638_ \atbs_core_0.spike_memory_0.n2406_o[18]\ _02634_ VPWR VGND _01901_ sg13g2_mux2_1
X_21833_ \atbs_core_0.spike_memory_0.n2362_o[18]\ \atbs_core_0.spike_memory_0.n2361_o[18]\ _02634_ VPWR VGND _01902_ sg13g2_mux2_1
X_21834_ \atbs_core_0.spike_memory_0.n2408_o[0]\ VPWR VGND _02639_ sg13g2_buf_1
X_21835_ _02639_ _02618_ _02634_ VPWR VGND _01903_ sg13g2_mux2_1
X_21836_ \atbs_core_0.spike_memory_0.n2408_o[1]\ VPWR VGND _02640_ sg13g2_buf_1
X_21837_ _02640_ _02619_ _02634_ VPWR VGND _01904_ sg13g2_mux2_1
X_21838_ \atbs_core_0.spike_memory_0.n2408_o[2]\ VPWR VGND _02641_ sg13g2_buf_1
X_21839_ _02641_ _02620_ _02634_ VPWR VGND _01905_ sg13g2_mux2_1
X_21840_ \atbs_core_0.spike_memory_0.n2408_o[3]\ VPWR VGND _02642_ sg13g2_buf_1
X_21841_ _02642_ _02621_ _02634_ VPWR VGND _01906_ sg13g2_mux2_1
X_21842_ \atbs_core_0.spike_memory_0.n2408_o[4]\ VPWR VGND _02643_ sg13g2_buf_1
X_21843_ _02613_ VPWR VGND _02644_ sg13g2_buf_1
X_21844_ _02643_ _02622_ _02644_ VPWR VGND _01907_ sg13g2_mux2_1
X_21845_ \atbs_core_0.spike_memory_0.n2408_o[5]\ VPWR VGND _02645_ sg13g2_buf_1
X_21846_ _02645_ _02623_ _02644_ VPWR VGND _01908_ sg13g2_mux2_1
X_21847_ \atbs_core_0.spike_memory_0.n2408_o[6]\ VPWR VGND _02646_ sg13g2_buf_1
X_21848_ _02646_ _02625_ _02644_ VPWR VGND _01909_ sg13g2_mux2_1
X_21849_ \atbs_core_0.spike_memory_0.n2408_o[7]\ VPWR VGND _02647_ sg13g2_buf_1
X_21850_ _02647_ _02626_ _02644_ VPWR VGND _01910_ sg13g2_mux2_1
X_21851_ \atbs_core_0.spike_memory_0.n2408_o[8]\ VPWR VGND _02648_ sg13g2_buf_1
X_21852_ _02648_ _02627_ _02644_ VPWR VGND _01911_ sg13g2_mux2_1
X_21853_ \atbs_core_0.spike_memory_0.n2408_o[9]\ VPWR VGND _02649_ sg13g2_buf_1
X_21854_ _02649_ _02628_ _02644_ VPWR VGND _01912_ sg13g2_mux2_1
X_21855_ _12625_ \atbs_core_0.spike_memory_0.n2362_o[0]\ _02644_ VPWR VGND _01913_ sg13g2_mux2_1
X_21856_ \atbs_core_0.spike_memory_0.n2408_o[10]\ VPWR VGND _02650_ sg13g2_buf_1
X_21857_ _02650_ _02629_ _02644_ VPWR VGND _01914_ sg13g2_mux2_1
X_21858_ \atbs_core_0.spike_memory_0.n2408_o[11]\ VPWR VGND _02651_ sg13g2_buf_1
X_21859_ _02651_ _02630_ _02644_ VPWR VGND _01915_ sg13g2_mux2_1
X_21860_ \atbs_core_0.spike_memory_0.n2408_o[12]\ VPWR VGND _02652_ sg13g2_buf_1
X_21861_ _02652_ _02631_ _02644_ VPWR VGND _01916_ sg13g2_mux2_1
X_21862_ \atbs_core_0.spike_memory_0.n2408_o[13]\ VPWR VGND _02653_ sg13g2_buf_1
X_21863_ _02191_ VPWR VGND _02654_ sg13g2_buf_1
X_21864_ _02653_ _02632_ _02654_ VPWR VGND _01917_ sg13g2_mux2_1
X_21865_ \atbs_core_0.spike_memory_0.n2408_o[14]\ VPWR VGND _02655_ sg13g2_buf_1
X_21866_ _02655_ _02633_ _02654_ VPWR VGND _01918_ sg13g2_mux2_1
X_21867_ \atbs_core_0.spike_memory_0.n2408_o[15]\ VPWR VGND _02656_ sg13g2_buf_1
X_21868_ _02656_ _02635_ _02654_ VPWR VGND _01919_ sg13g2_mux2_1
X_21869_ \atbs_core_0.spike_memory_0.n2408_o[16]\ VPWR VGND _02657_ sg13g2_buf_1
X_21870_ _02657_ _02636_ _02654_ VPWR VGND _01920_ sg13g2_mux2_1
X_21871_ \atbs_core_0.spike_memory_0.n2408_o[17]\ VPWR VGND _02658_ sg13g2_buf_1
X_21872_ _02658_ _02637_ _02654_ VPWR VGND _01921_ sg13g2_mux2_1
X_21873_ \atbs_core_0.spike_memory_0.n2408_o[18]\ VPWR VGND _02659_ sg13g2_buf_1
X_21874_ _02659_ _02638_ _02654_ VPWR VGND _01922_ sg13g2_mux2_1
X_21875_ \atbs_core_0.spike_memory_0.n2409_o[0]\ VPWR VGND _02660_ sg13g2_inv_1
X_21876_ _02639_ _02464_ VPWR VGND _02661_ sg13g2_nand2_1
X_21877_ _02660_ _02455_ _02661_ VPWR VGND _01923_ sg13g2_o21ai_1
X_21878_ _12630_ \atbs_core_0.spike_memory_0.n2362_o[1]\ _02654_ VPWR VGND _01924_ sg13g2_mux2_1
X_21879_ \atbs_core_0.spike_memory_0.n2409_o[1]\ VPWR VGND _02662_ sg13g2_inv_1
X_21880_ _02640_ _02464_ VPWR VGND _02663_ sg13g2_nand2_1
X_21881_ _02662_ _02455_ _02663_ VPWR VGND _01925_ sg13g2_o21ai_1
X_21882_ \atbs_core_0.spike_memory_0.n2409_o[2]\ VPWR VGND _02664_ sg13g2_inv_1
X_21883_ _12513_ VPWR VGND _02665_ sg13g2_buf_1
X_21884_ _02641_ _02464_ VPWR VGND _02666_ sg13g2_nand2_1
X_21885_ _02664_ _02665_ _02666_ VPWR VGND _01926_ sg13g2_o21ai_1
X_21886_ \atbs_core_0.spike_memory_0.n2409_o[3]\ VPWR VGND _02667_ sg13g2_inv_1
X_21887_ _02642_ _02464_ VPWR VGND _02668_ sg13g2_nand2_1
X_21888_ _02667_ _02665_ _02668_ VPWR VGND _01927_ sg13g2_o21ai_1
X_21889_ \atbs_core_0.spike_memory_0.n2409_o[4]\ VPWR VGND _02669_ sg13g2_inv_1
X_21890_ _02643_ _02464_ VPWR VGND _02670_ sg13g2_nand2_1
X_21891_ _02669_ _02665_ _02670_ VPWR VGND _01928_ sg13g2_o21ai_1
X_21892_ \atbs_core_0.spike_memory_0.n2409_o[5]\ _02645_ _02654_ VPWR VGND _01929_ sg13g2_mux2_1
X_21893_ \atbs_core_0.spike_memory_0.n2409_o[6]\ VPWR VGND _02671_ sg13g2_inv_1
X_21894_ _02646_ _02464_ VPWR VGND _02672_ sg13g2_nand2_1
X_21895_ _02671_ _02665_ _02672_ VPWR VGND _01930_ sg13g2_o21ai_1
X_21896_ \atbs_core_0.spike_memory_0.n2409_o[7]\ VPWR VGND _02673_ sg13g2_inv_1
X_21897_ _02191_ VPWR VGND _02674_ sg13g2_buf_1
X_21898_ _02647_ _02674_ VPWR VGND _02675_ sg13g2_nand2_1
X_21899_ _02673_ _02665_ _02675_ VPWR VGND _01931_ sg13g2_o21ai_1
X_21900_ \atbs_core_0.spike_memory_0.n2409_o[8]\ VPWR VGND _02676_ sg13g2_inv_1
X_21901_ _02648_ _02674_ VPWR VGND _02677_ sg13g2_nand2_1
X_21902_ _02676_ _02665_ _02677_ VPWR VGND _01932_ sg13g2_o21ai_1
X_21903_ \atbs_core_0.spike_memory_0.n2409_o[9]\ VPWR VGND _02678_ sg13g2_inv_1
X_21904_ _02649_ _02674_ VPWR VGND _02679_ sg13g2_nand2_1
X_21905_ _02678_ _02665_ _02679_ VPWR VGND _01933_ sg13g2_o21ai_1
X_21906_ \atbs_core_0.spike_memory_0.n2409_o[10]\ VPWR VGND _02680_ sg13g2_inv_1
X_21907_ _02650_ _02674_ VPWR VGND _02681_ sg13g2_nand2_1
X_21908_ _02680_ _02665_ _02681_ VPWR VGND _01934_ sg13g2_o21ai_1
X_21909_ _12643_ \atbs_core_0.spike_memory_0.n2362_o[2]\ _02654_ VPWR VGND _01935_ sg13g2_mux2_1
X_21910_ \atbs_core_0.spike_memory_0.n2409_o[11]\ _02651_ _02654_ VPWR VGND _01936_ sg13g2_mux2_1
X_21911_ \atbs_core_0.spike_memory_0.n2409_o[12]\ VPWR VGND _02682_ sg13g2_inv_1
X_21912_ _02652_ _02674_ VPWR VGND _02683_ sg13g2_nand2_1
X_21913_ _02682_ _02665_ _02683_ VPWR VGND _01937_ sg13g2_o21ai_1
X_21914_ _02191_ VPWR VGND _02684_ sg13g2_buf_1
X_21915_ \atbs_core_0.spike_memory_0.n2409_o[13]\ _02653_ _02684_ VPWR VGND _01938_ sg13g2_mux2_1
X_21916_ \atbs_core_0.spike_memory_0.n2409_o[14]\ VPWR VGND _02685_ sg13g2_inv_1
X_21917_ _02655_ _02674_ VPWR VGND _02686_ sg13g2_nand2_1
X_21918_ _02685_ _02665_ _02686_ VPWR VGND _01939_ sg13g2_o21ai_1
X_21919_ \atbs_core_0.spike_memory_0.n2409_o[15]\ VPWR VGND _02687_ sg13g2_inv_1
X_21920_ _02656_ _02674_ VPWR VGND _02688_ sg13g2_nand2_1
X_21921_ _02687_ _12514_ _02688_ VPWR VGND _01940_ sg13g2_o21ai_1
X_21922_ \atbs_core_0.spike_memory_0.n2409_o[16]\ VPWR VGND _02689_ sg13g2_inv_1
X_21923_ _02657_ _02674_ VPWR VGND _02690_ sg13g2_nand2_1
X_21924_ _02689_ _12514_ _02690_ VPWR VGND _01941_ sg13g2_o21ai_1
X_21925_ \atbs_core_0.spike_memory_0.n2409_o[17]\ VPWR VGND _02691_ sg13g2_inv_1
X_21926_ _02658_ _02674_ VPWR VGND _02692_ sg13g2_nand2_1
X_21927_ _02691_ _12514_ _02692_ VPWR VGND _01942_ sg13g2_o21ai_1
X_21928_ \atbs_core_0.spike_memory_0.n2409_o[18]\ VPWR VGND _02693_ sg13g2_inv_1
X_21929_ _02659_ _02674_ VPWR VGND _02694_ sg13g2_nand2_1
X_21930_ _02693_ _12514_ _02694_ VPWR VGND _01943_ sg13g2_o21ai_1
X_21931_ \atbs_core_0.spike_memory_0.n2410_o[0]\ \atbs_core_0.spike_memory_0.n2409_o[0]\ _02684_ VPWR VGND _01944_ sg13g2_mux2_1
X_21932_ \atbs_core_0.spike_memory_0.n2410_o[1]\ \atbs_core_0.spike_memory_0.n2409_o[1]\ _02684_ VPWR VGND _01945_ sg13g2_mux2_1
X_21933_ _12656_ \atbs_core_0.spike_memory_0.n2362_o[3]\ _02684_ VPWR VGND _01946_ sg13g2_mux2_1
X_21934_ \atbs_core_0.spike_memory_0.n2410_o[2]\ \atbs_core_0.spike_memory_0.n2409_o[2]\ _02684_ VPWR VGND _01947_ sg13g2_mux2_1
X_21935_ \atbs_core_0.spike_memory_0.n2410_o[3]\ \atbs_core_0.spike_memory_0.n2409_o[3]\ _02684_ VPWR VGND _01948_ sg13g2_mux2_1
X_21936_ \atbs_core_0.spike_memory_0.n2410_o[4]\ \atbs_core_0.spike_memory_0.n2409_o[4]\ _02684_ VPWR VGND _01949_ sg13g2_mux2_1
X_21937_ \atbs_core_0.spike_memory_0.n2410_o[5]\ \atbs_core_0.spike_memory_0.n2409_o[5]\ _02684_ VPWR VGND _01950_ sg13g2_mux2_1
X_21938_ \atbs_core_0.spike_memory_0.n2410_o[6]\ \atbs_core_0.spike_memory_0.n2409_o[6]\ _02684_ VPWR VGND _01951_ sg13g2_mux2_1
X_21939_ \atbs_core_0.spike_memory_0.n2410_o[7]\ \atbs_core_0.spike_memory_0.n2409_o[7]\ _02684_ VPWR VGND _01952_ sg13g2_mux2_1
X_21940_ \atbs_core_0.spike_memory_0.n2410_o[8]\ \atbs_core_0.spike_memory_0.n2409_o[8]\ _02182_ VPWR VGND _01953_ sg13g2_mux2_1
X_21941_ \atbs_core_0.spike_memory_0.n2410_o[9]\ \atbs_core_0.spike_memory_0.n2409_o[9]\ _02182_ VPWR VGND _01954_ sg13g2_mux2_1
X_21942_ \atbs_core_0.spike_memory_0.n2410_o[10]\ \atbs_core_0.spike_memory_0.n2409_o[10]\ _02182_ VPWR VGND _01955_ sg13g2_mux2_1
X_21943_ \atbs_core_0.spike_memory_0.n2410_o[11]\ \atbs_core_0.spike_memory_0.n2409_o[11]\ _02182_ VPWR VGND _01956_ sg13g2_mux2_1
X_21944_ _12669_ \atbs_core_0.spike_memory_0.n2362_o[4]\ _02182_ VPWR VGND _01957_ sg13g2_mux2_1
X_21945_ \atbs_core_0.spike_memory_0.n2358_o[9]\ \atbs_core_0.spike_memory_0.a_data[9]\ _02182_ VPWR VGND _01958_ sg13g2_mux2_1
X_21946_ \atbs_core_0.encoded_spike_strb\ \atbs_core_0.n1389_q\ VPWR VGND _02695_ sg13g2_nand2_1
X_21947_ _12248_ _02695_ VPWR VGND _02696_ sg13g2_nor2_1
X_21948_ _02696_ VPWR VGND _02697_ sg13g2_buf_1
X_21949_ _02697_ VPWR VGND \atbs_core_0.spike_memory_0.n2304_o\ sg13g2_buf_1
X_21950_ _07525_ VPWR VGND _02698_ sg13g2_buf_1
X_21951_ _02698_ VPWR VGND _02699_ sg13g2_buf_1
X_21952_ _02699_ VPWR VGND _02700_ sg13g2_buf_1
X_21953_ _02700_ VPWR VGND _02701_ sg13g2_buf_1
X_21954_ _02701_ VPWR VGND _02702_ sg13g2_buf_1
X_21955_ _02702_ \atbs_core_0.spike_memory_0.n2306_o[0]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01959_ sg13g2_mux2_1
X_21956_ _02702_ _02697_ VPWR VGND _02703_ sg13g2_nand2_1
X_21957_ _07523_ _02703_ VPWR VGND _01960_ sg13g2_xnor2_1
X_21958_ _02702_ _07523_ _02697_ VPWR VGND _02704_ sg13g2_nand3_1
X_21959_ _07520_ _02704_ VPWR VGND _01961_ sg13g2_xnor2_1
X_21960_ _02702_ _07523_ _07520_ _02697_ VPWR VGND 
+ _02705_
+ sg13g2_and4_1
X_21961_ _02705_ VPWR VGND _02706_ sg13g2_buf_1
X_21962_ _07517_ _02706_ VPWR VGND _01962_ sg13g2_xor2_1
X_21963_ _07517_ _02706_ VPWR VGND _02707_ sg13g2_nand2_1
X_21964_ _07537_ _02707_ VPWR VGND _01963_ sg13g2_xnor2_1
X_21965_ _07517_ _07537_ _02706_ VPWR VGND _02708_ sg13g2_nand3_1
X_21966_ \atbs_core_0.spike_memory_0.head[5]\ _02708_ VPWR VGND _01964_ sg13g2_xnor2_1
X_21967_ _07526_ VPWR VGND _02709_ sg13g2_buf_1
X_21968_ _02709_ VPWR VGND _02710_ sg13g2_buf_1
X_21969_ _02710_ VPWR VGND _02711_ sg13g2_buf_1
X_21970_ _02711_ VPWR VGND _02712_ sg13g2_buf_1
X_21971_ _02712_ VPWR VGND _02713_ sg13g2_buf_1
X_21972_ _02713_ VPWR VGND _02714_ sg13g2_buf_1
X_21973_ _02714_ \atbs_core_0.spike_memory_0.n2321_o[0]\ \atbs_core_0.spike_memory_0.n2319_o\ VPWR VGND _01965_ sg13g2_mux2_1
X_21974_ _02714_ \atbs_core_0.spike_memory_0.n2319_o\ VPWR VGND _02715_ sg13g2_nand2_1
X_21975_ _07522_ _02715_ VPWR VGND _01966_ sg13g2_xnor2_1
X_21976_ _02714_ _07522_ \atbs_core_0.spike_memory_0.n2319_o\ VPWR VGND _02716_ sg13g2_nand3_1
X_21977_ _07519_ _02716_ VPWR VGND _01967_ sg13g2_xnor2_1
X_21978_ _02714_ _07522_ _07519_ \atbs_core_0.spike_memory_0.n2319_o\ VPWR VGND 
+ _02717_
+ sg13g2_and4_1
X_21979_ _02717_ VPWR VGND _02718_ sg13g2_buf_1
X_21980_ _07518_ _02718_ VPWR VGND _01968_ sg13g2_xor2_1
X_21981_ _07518_ _02718_ VPWR VGND _02719_ sg13g2_nand2_1
X_21982_ _07538_ _02719_ VPWR VGND _01969_ sg13g2_xnor2_1
X_21983_ _07518_ _07538_ _02718_ VPWR VGND _02720_ sg13g2_nand3_1
X_21984_ \atbs_core_0.spike_memory_0.n2438_q[5]\ _02720_ VPWR VGND _01970_ sg13g2_xnor2_1
X_21985_ \atbs_core_0.spike_memory_0.a_data[0]\ \atbs_core_0.encoded_spike[0]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01971_ sg13g2_mux2_1
X_21986_ \atbs_core_0.spike_memory_0.a_data[10]\ \atbs_core_0.encoded_spike[10]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01972_ sg13g2_mux2_1
X_21987_ \atbs_core_0.spike_memory_0.a_data[11]\ \atbs_core_0.encoded_spike[11]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01973_ sg13g2_mux2_1
X_21988_ \atbs_core_0.spike_memory_0.a_data[12]\ \atbs_core_0.encoded_spike[12]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01974_ sg13g2_mux2_1
X_21989_ \atbs_core_0.spike_memory_0.a_data[13]\ \atbs_core_0.encoded_spike[13]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01975_ sg13g2_mux2_1
X_21990_ \atbs_core_0.spike_memory_0.a_data[14]\ \atbs_core_0.encoded_spike[14]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01976_ sg13g2_mux2_1
X_21991_ \atbs_core_0.spike_memory_0.a_data[15]\ \atbs_core_0.encoded_spike[15]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01977_ sg13g2_mux2_1
X_21992_ \atbs_core_0.spike_memory_0.a_data[16]\ \atbs_core_0.encoded_spike[16]\ \atbs_core_0.spike_memory_0.n2304_o\ VPWR VGND _01978_ sg13g2_mux2_1
X_21993_ _02697_ VPWR VGND _02721_ sg13g2_buf_1
X_21994_ \atbs_core_0.spike_memory_0.a_data[17]\ \atbs_core_0.encoded_spike[17]\ _02721_ VPWR VGND _01979_ sg13g2_mux2_1
X_21995_ \atbs_core_0.spike_memory_0.a_data[18]\ \atbs_core_0.encoded_spike[18]\ _02721_ VPWR VGND _01980_ sg13g2_mux2_1
X_21996_ \atbs_core_0.spike_memory_0.a_data[1]\ \atbs_core_0.encoded_spike[1]\ _02721_ VPWR VGND _01981_ sg13g2_mux2_1
X_21997_ \atbs_core_0.spike_memory_0.a_data[2]\ \atbs_core_0.encoded_spike[2]\ _02721_ VPWR VGND _01982_ sg13g2_mux2_1
X_21998_ \atbs_core_0.spike_memory_0.a_data[3]\ \atbs_core_0.encoded_spike[3]\ _02721_ VPWR VGND _01983_ sg13g2_mux2_1
X_21999_ \atbs_core_0.spike_memory_0.a_data[4]\ \atbs_core_0.encoded_spike[4]\ _02721_ VPWR VGND _01984_ sg13g2_mux2_1
X_22000_ \atbs_core_0.spike_memory_0.a_data[5]\ \atbs_core_0.encoded_spike[5]\ _02721_ VPWR VGND _01985_ sg13g2_mux2_1
X_22001_ \atbs_core_0.spike_memory_0.a_data[6]\ \atbs_core_0.encoded_spike[6]\ _02721_ VPWR VGND _01986_ sg13g2_mux2_1
X_22002_ \atbs_core_0.spike_memory_0.a_data[7]\ \atbs_core_0.encoded_spike[7]\ _02721_ VPWR VGND _01987_ sg13g2_mux2_1
X_22003_ \atbs_core_0.spike_memory_0.a_data[8]\ \atbs_core_0.encoded_spike[8]\ _02721_ VPWR VGND _01988_ sg13g2_mux2_1
X_22004_ \atbs_core_0.spike_memory_0.a_data[9]\ \atbs_core_0.encoded_spike[9]\ _02697_ VPWR VGND _01989_ sg13g2_mux2_1
X_22005_ _12017_ \atbs_core_0.spike_memory_0.n2319_o\ VPWR VGND _02722_ sg13g2_nor2_1
X_22006_ \atbs_core_0.spike_memory_0.n2333_o[0]\ \atbs_core_0.spike_memory_0.n2331_o\ _02722_ VPWR VGND _01990_ sg13g2_mux2_1
X_22007_ \atbs_core_0.spike_memory_0.n2331_o\ VPWR VGND _02723_ sg13g2_inv_1
X_22008_ \atbs_core_0.spike_memory_0.n2330_o\ \atbs_core_0.spike_memory_0.n2319_o\ _12018_ VPWR VGND _02724_ sg13g2_o21ai_1
X_22009_ _12018_ _02723_ _02724_ VPWR VGND _01991_ sg13g2_o21ai_1
X_22010_ \atbs_core_0.spike_memory_0.n2330_o\ VPWR VGND _02725_ sg13g2_inv_1
X_22011_ \atbs_core_0.spike_memory_0.n2317_o\ \atbs_core_0.spike_memory_0.n2319_o\ _12018_ VPWR VGND _02726_ sg13g2_o21ai_1
X_22012_ _12018_ _02725_ _02726_ VPWR VGND _01992_ sg13g2_o21ai_1
X_22013_ _07608_ VPWR VGND _02727_ sg13g2_inv_1
X_22014_ _07605_ _07601_ VPWR VGND _02728_ sg13g2_xor2_1
X_22015_ _02727_ _02728_ VPWR VGND _01993_ sg13g2_nor2_1
X_22016_ _07602_ _07607_ VPWR VGND _02729_ sg13g2_xor2_1
X_22017_ _02727_ _02729_ VPWR VGND _01994_ sg13g2_nor2_1
X_22018_ _07602_ _07605_ _07606_ VPWR VGND _02730_ sg13g2_nand3_1
X_22019_ _07603_ _02730_ VPWR VGND _02731_ sg13g2_xnor2_1
X_22020_ _07608_ _02731_ VPWR VGND _01995_ sg13g2_and2_1
X_22021_ _07602_ _07605_ VPWR VGND _02732_ sg13g2_nor2_1
X_22022_ _07603_ _02732_ VPWR VGND _02733_ sg13g2_nand2b_1
X_22023_ _07665_ _07668_ _07672_ VPWR VGND _02734_ sg13g2_nand3b_1
X_22024_ _07567_ _07675_ _07660_ _02727_ VPWR VGND 
+ _02735_
+ sg13g2_nor4_1
X_22025_ _02735_ VPWR VGND _02736_ sg13g2_inv_1
X_22026_ _02734_ _02736_ VPWR VGND _02737_ sg13g2_nor2_1
X_22027_ _02737_ VPWR VGND _02738_ sg13g2_buf_1
X_22028_ _07660_ _02727_ VPWR VGND _02739_ sg13g2_nor2_1
X_22029_ _07608_ _07660_ VPWR VGND _02740_ sg13g2_nor2b_1
X_22030_ _07673_ _02739_ _02740_ VPWR VGND _02741_ sg13g2_a21oi_1
X_22031_ _07660_ _02727_ _07675_ VPWR VGND _02742_ sg13g2_nand3b_1
X_22032_ _07675_ _02741_ _02742_ VPWR VGND _02743_ sg13g2_o21ai_1
X_22033_ _07568_ _07675_ _07660_ _07608_ VPWR VGND 
+ _02744_
+ sg13g2_nor4_1
X_22034_ _07568_ _02743_ _02744_ VPWR VGND _02745_ sg13g2_a21o_1
X_22035_ _02745_ VPWR VGND _02746_ sg13g2_buf_1
X_22036_ _02733_ _02738_ _02746_ VPWR VGND _02747_ sg13g2_a21oi_1
X_22037_ _07676_ _02736_ VPWR VGND _02748_ sg13g2_nor2_1
X_22038_ _02748_ VPWR VGND _02749_ sg13g2_buf_1
X_22039_ _02749_ _02747_ VPWR VGND _02750_ sg13g2_nand2_1
X_22040_ _07895_ _02747_ _02750_ VPWR VGND _01996_ sg13g2_o21ai_1
X_22041_ _07602_ _00063_ VPWR VGND _02751_ sg13g2_nor2_1
X_22042_ _07603_ _02751_ VPWR VGND _02752_ sg13g2_nand2b_1
X_22043_ _02738_ _02752_ _02746_ VPWR VGND _02753_ sg13g2_a21oi_1
X_22044_ _07880_ _02749_ _02753_ VPWR VGND _01997_ sg13g2_mux2_1
X_22045_ _07603_ _07602_ VPWR VGND _02754_ sg13g2_nor2b_1
X_22046_ _07605_ _02754_ VPWR VGND _02755_ sg13g2_nand2b_1
X_22047_ _02738_ _02755_ _02746_ VPWR VGND _02756_ sg13g2_a21oi_1
X_22048_ _07881_ _02749_ _02756_ VPWR VGND _01998_ sg13g2_mux2_1
X_22049_ _07605_ _02749_ _02754_ VPWR VGND _02757_ sg13g2_nand3_1
X_22050_ _07605_ _02754_ _02736_ VPWR VGND _02758_ sg13g2_a21oi_1
X_22051_ _02746_ _02758_ _07882_ VPWR VGND _02759_ sg13g2_o21ai_1
X_22052_ _02746_ _02757_ _02759_ VPWR VGND _01999_ sg13g2_o21ai_1
X_22053_ _07603_ _02732_ VPWR VGND _02760_ sg13g2_nand2_1
X_22054_ _02738_ _02760_ _02746_ VPWR VGND _02761_ sg13g2_a21oi_1
X_22055_ _02749_ _02761_ VPWR VGND _02762_ sg13g2_nand2_1
X_22056_ _07873_ _02761_ _02762_ VPWR VGND _02000_ sg13g2_o21ai_1
X_22057_ _07603_ _02751_ VPWR VGND _02763_ sg13g2_nand2_1
X_22058_ _02738_ _02763_ _02746_ VPWR VGND _02764_ sg13g2_a21oi_1
X_22059_ _07871_ _02749_ _02764_ VPWR VGND _02001_ sg13g2_mux2_1
X_22060_ _07605_ _07604_ _02738_ VPWR VGND _02765_ sg13g2_o21ai_1
X_22061_ _02746_ _02765_ VPWR VGND _02766_ sg13g2_nor2b_1
X_22062_ \atbs_core_0.uart_0.uart_rx_0.n3484_o\ _02749_ _02766_ VPWR VGND _02002_ sg13g2_mux2_1
X_22063_ _00063_ _07604_ _02738_ VPWR VGND _02767_ sg13g2_o21ai_1
X_22064_ _02746_ _02767_ VPWR VGND _02768_ sg13g2_nor2b_1
X_22065_ \atbs_core_0.uart_0.uart_rx_0.n3486_o\ _02749_ _02768_ VPWR VGND _02003_ sg13g2_mux2_1
X_22066_ _07644_ _07637_ VPWR VGND _02769_ sg13g2_xnor2_1
X_22067_ _07845_ _02769_ VPWR VGND _02004_ sg13g2_nor2_1
X_22068_ _07644_ _07637_ VPWR VGND _02770_ sg13g2_nand2_1
X_22069_ _07643_ _02770_ VPWR VGND _02771_ sg13g2_xor2_1
X_22070_ _07845_ _02771_ VPWR VGND _02005_ sg13g2_nor2_1
X_22071_ _00109_ _07847_ VPWR VGND _02772_ sg13g2_xnor2_1
X_22072_ _07846_ _02772_ _07637_ VPWR VGND _02773_ sg13g2_mux2_1
X_22073_ _07845_ _02773_ VPWR VGND _02006_ sg13g2_nor2_1
X_22074_ _07932_ VPWR VGND _02774_ sg13g2_buf_1
X_22075_ _08894_ _08495_ _02774_ VPWR VGND _00223_ sg13g2_mux2_1
X_22076_ _11159_ _08768_ _02774_ VPWR VGND _00224_ sg13g2_mux2_1
X_22077_ _07801_ VPWR VGND _02775_ sg13g2_buf_1
X_22078_ _02775_ VPWR VGND _02776_ sg13g2_buf_1
X_22079_ _08784_ _02776_ VPWR VGND _02777_ sg13g2_nand2_1
X_22080_ _11169_ _11321_ _02777_ VPWR VGND _00225_ sg13g2_o21ai_1
X_22081_ _11141_ _11343_ VPWR VGND _02778_ sg13g2_nand2_1
X_22082_ _08767_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02778_ VPWR VGND _00226_ sg13g2_o21ai_1
X_22083_ _11140_ _08765_ _02774_ VPWR VGND _00227_ sg13g2_mux2_1
X_22084_ _11143_ _08795_ _02774_ VPWR VGND _00228_ sg13g2_mux2_1
X_22085_ _11180_ _08794_ _02774_ VPWR VGND _00229_ sg13g2_mux2_1
X_22086_ _11138_ _11343_ VPWR VGND _02779_ sg13g2_nand2_1
X_22087_ _08764_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02779_ VPWR VGND _00230_ sg13g2_o21ai_1
X_22088_ _11187_ _11343_ VPWR VGND _02780_ sg13g2_nand2_1
X_22089_ _08819_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02780_ VPWR VGND _00231_ sg13g2_o21ai_1
X_22090_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ _11335_ VPWR VGND _00232_ sg13g2_mux2_1
X_22091_ _09070_ _08890_ _11335_ VPWR VGND _00233_ sg13g2_mux2_1
X_22092_ _08435_ _02776_ VPWR VGND _02781_ sg13g2_nand2_1
X_22093_ _08860_ _11321_ _02781_ VPWR VGND _00234_ sg13g2_o21ai_1
X_22094_ _08977_ VPWR VGND _02782_ sg13g2_buf_1
X_22095_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _02776_ VPWR VGND _02783_ sg13g2_nand2_1
X_22096_ _08887_ _02782_ _02783_ VPWR VGND _00235_ sg13g2_o21ai_1
X_22097_ _09064_ _02776_ VPWR VGND _02784_ sg13g2_nand2_1
X_22098_ _08886_ _02782_ _02784_ VPWR VGND _00236_ sg13g2_o21ai_1
X_22099_ _10285_ VPWR VGND _02785_ sg13g2_buf_1
X_22100_ _09065_ _02785_ VPWR VGND _02786_ sg13g2_nand2_1
X_22101_ _08881_ _02782_ _02786_ VPWR VGND _00237_ sg13g2_o21ai_1
X_22102_ _09062_ _02785_ VPWR VGND _02787_ sg13g2_nand2_1
X_22103_ _08880_ _02782_ _02787_ VPWR VGND _00238_ sg13g2_o21ai_1
X_22104_ _09000_ _08771_ _11335_ VPWR VGND _00239_ sg13g2_mux2_1
X_22105_ _09001_ _08772_ _11335_ VPWR VGND _00240_ sg13g2_mux2_1
X_22106_ _08998_ _08769_ _11335_ VPWR VGND _00241_ sg13g2_mux2_1
X_22107_ _08996_ _02785_ VPWR VGND _02788_ sg13g2_nand2_1
X_22108_ _08777_ _02782_ _02788_ VPWR VGND _00242_ sg13g2_o21ai_1
X_22109_ _08990_ _08768_ _11335_ VPWR VGND _00243_ sg13g2_mux2_1
X_22110_ _08987_ _08784_ _11335_ VPWR VGND _00244_ sg13g2_mux2_1
X_22111_ _12415_ _11343_ VPWR VGND _02789_ sg13g2_nand2_1
X_22112_ _08410_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02789_ VPWR VGND _00245_ sg13g2_o21ai_1
X_22113_ _08988_ _02785_ VPWR VGND _02790_ sg13g2_nand2_1
X_22114_ _08767_ _02782_ _02790_ VPWR VGND _00246_ sg13g2_o21ai_1
X_22115_ _08986_ _08765_ _11335_ VPWR VGND _00247_ sg13g2_mux2_1
X_22116_ _09016_ _08795_ _11335_ VPWR VGND _00248_ sg13g2_mux2_1
X_22117_ _08970_ VPWR VGND _02791_ sg13g2_buf_1
X_22118_ _08985_ _08794_ _02791_ VPWR VGND _00249_ sg13g2_mux2_1
X_22119_ _08983_ _02785_ VPWR VGND _02792_ sg13g2_nand2_1
X_22120_ _08764_ _02782_ _02792_ VPWR VGND _00250_ sg13g2_o21ai_1
X_22121_ _09031_ _02785_ VPWR VGND _02793_ sg13g2_nand2_1
X_22122_ _08819_ _02782_ _02793_ VPWR VGND _00251_ sg13g2_o21ai_1
X_22123_ _07932_ VPWR VGND _02794_ sg13g2_buf_1
X_22124_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ _02794_ VPWR VGND _00252_ sg13g2_mux2_1
X_22125_ _09070_ _09242_ _02794_ VPWR VGND _00253_ sg13g2_mux2_1
X_22126_ _09240_ _02785_ VPWR VGND _02795_ sg13g2_nand2_1
X_22127_ _09069_ _02782_ _02795_ VPWR VGND _00254_ sg13g2_o21ai_1
X_22128_ _09064_ _11343_ VPWR VGND _02796_ sg13g2_nand2_1
X_22129_ _09238_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02796_ VPWR VGND _00255_ sg13g2_o21ai_1
X_22130_ _08457_ _02785_ VPWR VGND _02797_ sg13g2_nand2_1
X_22131_ _08569_ _02782_ _02797_ VPWR VGND _00256_ sg13g2_o21ai_1
X_22132_ _09065_ _11343_ VPWR VGND _02798_ sg13g2_nand2_1
X_22133_ _09239_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02798_ VPWR VGND _00257_ sg13g2_o21ai_1
X_22134_ _09062_ _09237_ _02794_ VPWR VGND _00258_ sg13g2_mux2_1
X_22135_ _09000_ _11343_ VPWR VGND _02799_ sg13g2_nand2_1
X_22136_ _09256_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ _02799_ VPWR VGND _00259_ sg13g2_o21ai_1
X_22137_ _09001_ _09176_ _02794_ VPWR VGND _00260_ sg13g2_mux2_1
X_22138_ _08998_ _09173_ _02794_ VPWR VGND _00261_ sg13g2_mux2_1
X_22139_ _07931_ VPWR VGND _02800_ sg13g2_buf_1
X_22140_ _02800_ VPWR VGND _02801_ sg13g2_buf_1
X_22141_ _09181_ _02785_ VPWR VGND _02802_ sg13g2_nand2_1
X_22142_ _08997_ _02801_ _02802_ VPWR VGND _00262_ sg13g2_o21ai_1
X_22143_ _08990_ _09168_ _02794_ VPWR VGND _00263_ sg13g2_mux2_1
X_22144_ _08987_ _09165_ _02794_ VPWR VGND _00264_ sg13g2_mux2_1
X_22145_ _08988_ _09166_ _02794_ VPWR VGND _00265_ sg13g2_mux2_1
X_22146_ _08981_ VPWR VGND _02803_ sg13g2_buf_1
X_22147_ _08986_ _11343_ VPWR VGND _02804_ sg13g2_nand2_1
X_22148_ _09198_ _02803_ _02804_ VPWR VGND _00266_ sg13g2_o21ai_1
X_22149_ _08465_ _02785_ VPWR VGND _02805_ sg13g2_nand2_1
X_22150_ _12443_ _02801_ _02805_ VPWR VGND _00267_ sg13g2_o21ai_1
X_22151_ _09016_ _09192_ _02794_ VPWR VGND _00268_ sg13g2_mux2_1
X_22152_ _08985_ _09163_ _02794_ VPWR VGND _00269_ sg13g2_mux2_1
X_22153_ _10285_ VPWR VGND _02806_ sg13g2_buf_1
X_22154_ _09162_ _02806_ VPWR VGND _02807_ sg13g2_nand2_1
X_22155_ _08984_ _02801_ _02807_ VPWR VGND _00270_ sg13g2_o21ai_1
X_22156_ _09155_ _02806_ VPWR VGND _02808_ sg13g2_nand2_1
X_22157_ _09143_ _02801_ _02808_ VPWR VGND _00271_ sg13g2_o21ai_1
X_22158_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ _02791_ VPWR VGND _00272_ sg13g2_mux2_1
X_22159_ _09466_ _09242_ _02791_ VPWR VGND _00273_ sg13g2_mux2_1
X_22160_ _09464_ _09240_ _02791_ VPWR VGND _00274_ sg13g2_mux2_1
X_22161_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ _02806_ VPWR VGND _02809_ sg13g2_nand2_1
X_22162_ _09238_ _02801_ _02809_ VPWR VGND _00275_ sg13g2_o21ai_1
X_22163_ _09462_ _02806_ VPWR VGND _02810_ sg13g2_nand2_1
X_22164_ _09239_ _02801_ _02810_ VPWR VGND _00276_ sg13g2_o21ai_1
X_22165_ _09483_ _09237_ _02791_ VPWR VGND _00277_ sg13g2_mux2_1
X_22166_ _08654_ _02806_ VPWR VGND _02811_ sg13g2_nand2_1
X_22167_ _09868_ _02801_ _02811_ VPWR VGND _00278_ sg13g2_o21ai_1
X_22168_ _09362_ _02806_ VPWR VGND _02812_ sg13g2_nand2_1
X_22169_ _09256_ _02801_ _02812_ VPWR VGND _00279_ sg13g2_o21ai_1
X_22170_ _09363_ _09176_ _02791_ VPWR VGND _00280_ sg13g2_mux2_1
X_22171_ _09357_ _09173_ _02791_ VPWR VGND _00281_ sg13g2_mux2_1
X_22172_ _09356_ _02806_ VPWR VGND _02813_ sg13g2_nand2_1
X_22173_ _09182_ _02801_ _02813_ VPWR VGND _00282_ sg13g2_o21ai_1
X_22174_ _09368_ _09168_ _02791_ VPWR VGND _00283_ sg13g2_mux2_1
X_22175_ _09165_ _11343_ VPWR VGND _02814_ sg13g2_nand2_1
X_22176_ _09355_ _02803_ _02814_ VPWR VGND _00284_ sg13g2_o21ai_1
X_22177_ _09352_ _09166_ _02791_ VPWR VGND _00285_ sg13g2_mux2_1
X_22178_ _09351_ _02806_ VPWR VGND _02815_ sg13g2_nand2_1
X_22179_ _09198_ _02801_ _02815_ VPWR VGND _00286_ sg13g2_o21ai_1
X_22180_ _09413_ _09192_ _02791_ VPWR VGND _00287_ sg13g2_mux2_1
X_22181_ _10628_ VPWR VGND _02816_ sg13g2_buf_1
X_22182_ _09163_ _02816_ VPWR VGND _02817_ sg13g2_nand2_1
X_22183_ _09401_ _02803_ _02817_ VPWR VGND _00288_ sg13g2_o21ai_1
X_22184_ _12449_ _02816_ VPWR VGND _02818_ sg13g2_nand2_1
X_22185_ _08694_ _02803_ _02818_ VPWR VGND _00289_ sg13g2_o21ai_1
X_22186_ _08970_ VPWR VGND _02819_ sg13g2_buf_1
X_22187_ _09347_ _09162_ _02819_ VPWR VGND _00290_ sg13g2_mux2_1
X_22188_ _09346_ VPWR VGND _02820_ sg13g2_inv_1
X_22189_ _09155_ _02816_ VPWR VGND _02821_ sg13g2_nand2_1
X_22190_ _02820_ _02803_ _02821_ VPWR VGND _00291_ sg13g2_o21ai_1
X_22191_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ _02819_ VPWR VGND _00292_ sg13g2_mux2_1
X_22192_ _09630_ _09466_ _02819_ VPWR VGND _00293_ sg13g2_mux2_1
X_22193_ _09628_ _09464_ _02819_ VPWR VGND _00294_ sg13g2_mux2_1
X_22194_ _02800_ VPWR VGND _02822_ sg13g2_buf_1
X_22195_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _02806_ VPWR VGND _02823_ sg13g2_nand2_1
X_22196_ _09471_ _02822_ _02823_ VPWR VGND _00295_ sg13g2_o21ai_1
X_22197_ _09626_ _09462_ _02819_ VPWR VGND _00296_ sg13g2_mux2_1
X_22198_ _09624_ _09483_ _02819_ VPWR VGND _00297_ sg13g2_mux2_1
X_22199_ _09555_ _09362_ _02819_ VPWR VGND _00298_ sg13g2_mux2_1
X_22200_ _09363_ _02816_ VPWR VGND _02824_ sg13g2_nand2_1
X_22201_ _09554_ _02803_ _02824_ VPWR VGND _00299_ sg13g2_o21ai_1
X_22202_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[16]\ _02806_ VPWR VGND _02825_ sg13g2_nand2_1
X_22203_ _09035_ _02822_ _02825_ VPWR VGND _00300_ sg13g2_o21ai_1
X_22204_ _09550_ _09357_ _02819_ VPWR VGND _00301_ sg13g2_mux2_1
X_22205_ _02775_ VPWR VGND _02826_ sg13g2_buf_1
X_22206_ _09549_ _02826_ VPWR VGND _02827_ sg13g2_nand2_1
X_22207_ _09373_ _02822_ _02827_ VPWR VGND _00302_ sg13g2_o21ai_1
X_22208_ _09560_ _09368_ _02819_ VPWR VGND _00303_ sg13g2_mux2_1
X_22209_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[11]\ _02826_ VPWR VGND _02828_ sg13g2_nand2_1
X_22210_ _09355_ _02822_ _02828_ VPWR VGND _00304_ sg13g2_o21ai_1
X_22211_ _09540_ _09352_ _02819_ VPWR VGND _00305_ sg13g2_mux2_1
X_22212_ _09546_ _02826_ VPWR VGND _02829_ sg13g2_nand2_1
X_22213_ _09433_ _02822_ _02829_ VPWR VGND _00306_ sg13g2_o21ai_1
X_22214_ _10628_ VPWR VGND _02830_ sg13g2_buf_1
X_22215_ _09542_ _09413_ _02830_ VPWR VGND _00307_ sg13g2_mux2_1
X_22216_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[15]\ _02826_ VPWR VGND _02831_ sg13g2_nand2_1
X_22217_ _09401_ _02822_ _02831_ VPWR VGND _00308_ sg13g2_o21ai_1
X_22218_ _09675_ _09347_ _02830_ VPWR VGND _00309_ sg13g2_mux2_1
X_22219_ _09684_ _02826_ VPWR VGND _02832_ sg13g2_nand2_1
X_22220_ _02820_ _02822_ _02832_ VPWR VGND _00310_ sg13g2_o21ai_1
X_22221_ _08713_ _02826_ VPWR VGND _02833_ sg13g2_nand2_1
X_22222_ _08762_ _02822_ _02833_ VPWR VGND _00311_ sg13g2_o21ai_1
X_22223_ _07932_ VPWR VGND _02834_ sg13g2_buf_1
X_22224_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ _02834_ VPWR VGND _00312_ sg13g2_mux2_1
X_22225_ _09630_ _09804_ _02834_ VPWR VGND _00313_ sg13g2_mux2_1
X_22226_ _09628_ _02816_ VPWR VGND _02835_ sg13g2_nand2_1
X_22227_ _09803_ _02803_ _02835_ VPWR VGND _00314_ sg13g2_o21ai_1
X_22228_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _02816_ VPWR VGND _02836_ sg13g2_nand2_1
X_22229_ _09802_ _02803_ _02836_ VPWR VGND _00315_ sg13g2_o21ai_1
X_22230_ _09626_ _09810_ _02834_ VPWR VGND _00316_ sg13g2_mux2_1
X_22231_ _09624_ _02816_ VPWR VGND _02837_ sg13g2_nand2_1
X_22232_ _09788_ _02803_ _02837_ VPWR VGND _00317_ sg13g2_o21ai_1
X_22233_ _09555_ _09730_ _02834_ VPWR VGND _00318_ sg13g2_mux2_1
X_22234_ _09731_ _02826_ VPWR VGND _02838_ sg13g2_nand2_1
X_22235_ _09554_ _02822_ _02838_ VPWR VGND _00319_ sg13g2_o21ai_1
X_22236_ _09550_ _09728_ _02834_ VPWR VGND _00320_ sg13g2_mux2_1
X_22237_ _09738_ _02826_ VPWR VGND _02839_ sg13g2_nand2_1
X_22238_ _09565_ _02822_ _02839_ VPWR VGND _00321_ sg13g2_o21ai_1
X_22239_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ _08495_ _02830_ VPWR VGND _00322_ sg13g2_mux2_1
X_22240_ _09560_ _09725_ _02834_ VPWR VGND _00323_ sg13g2_mux2_1
X_22241_ _02800_ VPWR VGND _02840_ sg13g2_buf_1
X_22242_ _09724_ _02826_ VPWR VGND _02841_ sg13g2_nand2_1
X_22243_ _09570_ _02840_ _02841_ VPWR VGND _00324_ sg13g2_o21ai_1
X_22244_ _09540_ _09748_ _02834_ VPWR VGND _00325_ sg13g2_mux2_1
X_22245_ _09546_ _09752_ _02834_ VPWR VGND _00326_ sg13g2_mux2_1
X_22246_ _09542_ _09717_ _02834_ VPWR VGND _00327_ sg13g2_mux2_1
X_22247_ _09715_ _02826_ VPWR VGND _02842_ sg13g2_nand2_1
X_22248_ _09676_ _02840_ _02842_ VPWR VGND _00328_ sg13g2_o21ai_1
X_22249_ _09675_ _09888_ _02834_ VPWR VGND _00329_ sg13g2_mux2_1
X_22250_ _07932_ VPWR VGND _02843_ sg13g2_buf_1
X_22251_ _09684_ _09896_ _02843_ VPWR VGND _00330_ sg13g2_mux2_1
X_22252_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ _02843_ VPWR VGND _00331_ sg13g2_mux2_1
X_22253_ _09804_ _10014_ _02843_ VPWR VGND _00332_ sg13g2_mux2_1
X_22254_ _10723_ _08497_ _02830_ VPWR VGND _00333_ sg13g2_mux2_1
X_22255_ _08892_ _08497_ _02843_ VPWR VGND _00334_ sg13g2_mux2_1
X_22256_ _02775_ VPWR VGND _02844_ sg13g2_buf_1
X_22257_ _10012_ _02844_ VPWR VGND _02845_ sg13g2_nand2_1
X_22258_ _09803_ _02840_ _02845_ VPWR VGND _00335_ sg13g2_o21ai_1
X_22259_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _02844_ VPWR VGND _02846_ sg13g2_nand2_1
X_22260_ _09802_ _02840_ _02846_ VPWR VGND _00336_ sg13g2_o21ai_1
X_22261_ _09810_ _02816_ VPWR VGND _02847_ sg13g2_nand2_1
X_22262_ _10011_ _02803_ _02847_ VPWR VGND _00337_ sg13g2_o21ai_1
X_22263_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ _02844_ VPWR VGND _02848_ sg13g2_nand2_1
X_22264_ _09788_ _02840_ _02848_ VPWR VGND _00338_ sg13g2_o21ai_1
X_22265_ _09730_ _09923_ _02843_ VPWR VGND _00339_ sg13g2_mux2_1
X_22266_ _09731_ _09924_ _02843_ VPWR VGND _00340_ sg13g2_mux2_1
X_22267_ _09728_ _09921_ _02843_ VPWR VGND _00341_ sg13g2_mux2_1
X_22268_ _09929_ _02844_ VPWR VGND _02849_ sg13g2_nand2_1
X_22269_ _09739_ _02840_ _02849_ VPWR VGND _00342_ sg13g2_o21ai_1
X_22270_ _08981_ VPWR VGND _02850_ sg13g2_buf_1
X_22271_ _09725_ _02816_ VPWR VGND _02851_ sg13g2_nand2_1
X_22272_ _09939_ _02850_ _02851_ VPWR VGND _00343_ sg13g2_o21ai_1
X_22273_ _09919_ _02844_ VPWR VGND _02852_ sg13g2_nand2_1
X_22274_ _09762_ _02840_ _02852_ VPWR VGND _00344_ sg13g2_o21ai_1
X_22275_ _08492_ _02816_ VPWR VGND _02853_ sg13g2_nand2_1
X_22276_ _10722_ _02850_ _02853_ VPWR VGND _00345_ sg13g2_o21ai_1
X_22277_ _10628_ VPWR VGND _02854_ sg13g2_buf_1
X_22278_ _09748_ _02854_ VPWR VGND _02855_ sg13g2_nand2_1
X_22279_ _09918_ _02850_ _02855_ VPWR VGND _00346_ sg13g2_o21ai_1
X_22280_ _09752_ _09943_ _02843_ VPWR VGND _00347_ sg13g2_mux2_1
X_22281_ _09717_ _02854_ VPWR VGND _02856_ sg13g2_nand2_1
X_22282_ _09964_ _02850_ _02856_ VPWR VGND _00348_ sg13g2_o21ai_1
X_22283_ _09715_ _09968_ _02843_ VPWR VGND _00349_ sg13g2_mux2_1
X_22284_ _09888_ _10076_ _02843_ VPWR VGND _00350_ sg13g2_mux2_1
X_22285_ _09896_ _02854_ VPWR VGND _02857_ sg13g2_nand2_1
X_22286_ _10097_ _02850_ _02857_ VPWR VGND _00351_ sg13g2_o21ai_1
X_22287_ _07932_ VPWR VGND _02858_ sg13g2_buf_1
X_22288_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ _02858_ VPWR VGND _00352_ sg13g2_mux2_1
X_22289_ _10014_ _10217_ _02858_ VPWR VGND _00353_ sg13g2_mux2_1
X_22290_ _10012_ _10221_ _02858_ VPWR VGND _00354_ sg13g2_mux2_1
X_22291_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ _02844_ VPWR VGND _02859_ sg13g2_nand2_1
X_22292_ _10010_ _02840_ _02859_ VPWR VGND _00355_ sg13g2_o21ai_1
X_22293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[22]\ _02844_ VPWR VGND _02860_ sg13g2_nand2_1
X_22294_ _08488_ _02840_ _02860_ VPWR VGND _00356_ sg13g2_o21ai_1
X_22295_ _10214_ _02844_ VPWR VGND _02861_ sg13g2_nand2_1
X_22296_ _10011_ _02840_ _02861_ VPWR VGND _00357_ sg13g2_o21ai_1
X_22297_ _02800_ VPWR VGND _02862_ sg13g2_buf_1
X_22298_ _10212_ _02844_ VPWR VGND _02863_ sg13g2_nand2_1
X_22299_ _10023_ _02862_ _02863_ VPWR VGND _00358_ sg13g2_o21ai_1
X_22300_ _09923_ _02854_ VPWR VGND _02864_ sg13g2_nand2_1
X_22301_ _10196_ _02850_ _02864_ VPWR VGND _00359_ sg13g2_o21ai_1
X_22302_ _09924_ _10128_ _02858_ VPWR VGND _00360_ sg13g2_mux2_1
X_22303_ _09921_ _02854_ VPWR VGND _02865_ sg13g2_nand2_1
X_22304_ _10126_ _02850_ _02865_ VPWR VGND _00361_ sg13g2_o21ai_1
X_22305_ _10123_ _02844_ VPWR VGND _02866_ sg13g2_nand2_1
X_22306_ _09930_ _02862_ _02866_ VPWR VGND _00362_ sg13g2_o21ai_1
X_22307_ _02775_ VPWR VGND _02867_ sg13g2_buf_1
X_22308_ _10121_ _02867_ VPWR VGND _02868_ sg13g2_nand2_1
X_22309_ _09939_ _02862_ _02868_ VPWR VGND _00363_ sg13g2_o21ai_1
X_22310_ _09919_ _10143_ _02858_ VPWR VGND _00364_ sg13g2_mux2_1
X_22311_ _10119_ _02867_ VPWR VGND _02869_ sg13g2_nand2_1
X_22312_ _09918_ _02862_ _02869_ VPWR VGND _00365_ sg13g2_o21ai_1
X_22313_ _09943_ _02854_ VPWR VGND _02870_ sg13g2_nand2_1
X_22314_ _10148_ _02850_ _02870_ VPWR VGND _00366_ sg13g2_o21ai_1
X_22315_ _10729_ _08483_ _02830_ VPWR VGND _00367_ sg13g2_mux2_1
X_22316_ _10153_ _02867_ VPWR VGND _02871_ sg13g2_nand2_1
X_22317_ _09964_ _02862_ _02871_ VPWR VGND _00368_ sg13g2_o21ai_1
X_22318_ _09968_ _10157_ _02858_ VPWR VGND _00369_ sg13g2_mux2_1
X_22319_ _10076_ _10117_ _02858_ VPWR VGND _00370_ sg13g2_mux2_1
X_22320_ _10164_ _02867_ VPWR VGND _02872_ sg13g2_nand2_1
X_22321_ _10097_ _02862_ _02872_ VPWR VGND _00371_ sg13g2_o21ai_1
X_22322_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ _02858_ VPWR VGND _00372_ sg13g2_mux2_1
X_22323_ _10217_ _10385_ _02858_ VPWR VGND _00373_ sg13g2_mux2_1
X_22324_ _10221_ _10383_ _02858_ VPWR VGND _00374_ sg13g2_mux2_1
X_22325_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ _02867_ VPWR VGND _02873_ sg13g2_nand2_1
X_22326_ _10216_ _02862_ _02873_ VPWR VGND _00375_ sg13g2_o21ai_1
X_22327_ _10285_ VPWR VGND _02874_ sg13g2_buf_1
X_22328_ _10214_ _10371_ _02874_ VPWR VGND _00376_ sg13g2_mux2_1
X_22329_ _10212_ _10370_ _02874_ VPWR VGND _00377_ sg13g2_mux2_1
X_22330_ _10736_ _08478_ _02830_ VPWR VGND _00378_ sg13g2_mux2_1
X_22331_ _10308_ _02867_ VPWR VGND _02875_ sg13g2_nand2_1
X_22332_ _10196_ _02862_ _02875_ VPWR VGND _00379_ sg13g2_o21ai_1
X_22333_ _10128_ _10309_ _02874_ VPWR VGND _00380_ sg13g2_mux2_1
X_22334_ _10306_ _02867_ VPWR VGND _02876_ sg13g2_nand2_1
X_22335_ _10126_ _02862_ _02876_ VPWR VGND _00381_ sg13g2_o21ai_1
X_22336_ _10305_ _02867_ VPWR VGND _02877_ sg13g2_nand2_1
X_22337_ _10133_ _02862_ _02877_ VPWR VGND _00382_ sg13g2_o21ai_1
X_22338_ _10121_ _10313_ _02874_ VPWR VGND _00383_ sg13g2_mux2_1
X_22339_ _10143_ _10304_ _02874_ VPWR VGND _00384_ sg13g2_mux2_1
X_22340_ _10119_ _10299_ _02874_ VPWR VGND _00385_ sg13g2_mux2_1
X_22341_ _02800_ VPWR VGND _02878_ sg13g2_buf_1
X_22342_ _10296_ _02867_ VPWR VGND _02879_ sg13g2_nand2_1
X_22343_ _10148_ _02878_ _02879_ VPWR VGND _00386_ sg13g2_o21ai_1
X_22344_ _10153_ _10297_ _02874_ VPWR VGND _00387_ sg13g2_mux2_1
X_22345_ _10157_ _10295_ _02874_ VPWR VGND _00388_ sg13g2_mux2_1
X_22346_ _10646_ _02867_ VPWR VGND _02880_ sg13g2_nand2_1
X_22347_ _08511_ _02878_ _02880_ VPWR VGND _00389_ sg13g2_o21ai_1
X_22348_ _10117_ _10293_ _02874_ VPWR VGND _00390_ sg13g2_mux2_1
X_22349_ _10164_ _10292_ _02874_ VPWR VGND _00391_ sg13g2_mux2_1
X_22350_ _10285_ VPWR VGND _02881_ sg13g2_buf_1
X_22351_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ _02881_ VPWR VGND _00392_ sg13g2_mux2_1
X_22352_ _10385_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ _02881_ VPWR VGND _00393_ sg13g2_mux2_1
X_22353_ _10383_ _02854_ VPWR VGND _02882_ sg13g2_nand2_1
X_22354_ _10556_ _02850_ _02882_ VPWR VGND _00394_ sg13g2_o21ai_1
X_22355_ _02775_ VPWR VGND _02883_ sg13g2_buf_1
X_22356_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ _02883_ VPWR VGND _02884_ sg13g2_nand2_1
X_22357_ _10382_ _02878_ _02884_ VPWR VGND _00395_ sg13g2_o21ai_1
X_22358_ _10371_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _02881_ VPWR VGND _00396_ sg13g2_mux2_1
X_22359_ _10370_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _02881_ VPWR VGND _00397_ sg13g2_mux2_1
X_22360_ _10473_ _02883_ VPWR VGND _02885_ sg13g2_nand2_1
X_22361_ _10377_ _02878_ _02885_ VPWR VGND _00398_ sg13g2_o21ai_1
X_22362_ _10309_ _10474_ _02881_ VPWR VGND _00399_ sg13g2_mux2_1
X_22363_ _10647_ _08428_ _02830_ VPWR VGND _00400_ sg13g2_mux2_1
X_22364_ _10306_ _02854_ VPWR VGND _02886_ sg13g2_nand2_1
X_22365_ _10472_ _02850_ _02886_ VPWR VGND _00401_ sg13g2_o21ai_1
X_22366_ _10470_ _02883_ VPWR VGND _02887_ sg13g2_nand2_1
X_22367_ _10318_ _02878_ _02887_ VPWR VGND _00402_ sg13g2_o21ai_1
X_22368_ _10313_ _10480_ _02881_ VPWR VGND _00403_ sg13g2_mux2_1
X_22369_ _10304_ _10487_ _02881_ VPWR VGND _00404_ sg13g2_mux2_1
X_22370_ _10299_ _10464_ _02881_ VPWR VGND _00405_ sg13g2_mux2_1
X_22371_ _10461_ _02883_ VPWR VGND _02888_ sg13g2_nand2_1
X_22372_ _10327_ _02878_ _02888_ VPWR VGND _00406_ sg13g2_o21ai_1
X_22373_ _10297_ _10462_ _02881_ VPWR VGND _00407_ sg13g2_mux2_1
X_22374_ _08970_ VPWR VGND _02889_ sg13g2_buf_1
X_22375_ _10295_ _02854_ VPWR VGND _02890_ sg13g2_nand2_1
X_22376_ _10460_ _02889_ _02890_ VPWR VGND _00408_ sg13g2_o21ai_1
X_22377_ _10293_ _10501_ _02881_ VPWR VGND _00409_ sg13g2_mux2_1
X_22378_ _10292_ _02854_ VPWR VGND _02891_ sg13g2_nand2_1
X_22379_ _10607_ _02889_ _02891_ VPWR VGND _00410_ sg13g2_o21ai_1
X_22380_ _10643_ _08418_ _02830_ VPWR VGND _00411_ sg13g2_mux2_1
X_22381_ _10642_ _02883_ VPWR VGND _02892_ sg13g2_nand2_1
X_22382_ _08444_ _02878_ _02892_ VPWR VGND _00412_ sg13g2_o21ai_1
X_22383_ _10652_ _08435_ _02830_ VPWR VGND _00413_ sg13g2_mux2_1
X_22384_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[11]\ _02883_ VPWR VGND _02893_ sg13g2_nand2_1
X_22385_ _08410_ _02878_ _02893_ VPWR VGND _00414_ sg13g2_o21ai_1
X_22386_ _08492_ _02883_ VPWR VGND _02894_ sg13g2_nand2_1
X_22387_ _08889_ _02878_ _02894_ VPWR VGND _00415_ sg13g2_o21ai_1
X_22388_ _10636_ _08457_ _02830_ VPWR VGND _00416_ sg13g2_mux2_1
X_22389_ _10635_ _02883_ VPWR VGND _02895_ sg13g2_nand2_1
X_22390_ _08663_ _02878_ _02895_ VPWR VGND _00417_ sg13g2_o21ai_1
X_22391_ _10628_ VPWR VGND _02896_ sg13g2_buf_1
X_22392_ _10676_ _08654_ _02896_ VPWR VGND _00418_ sg13g2_mux2_1
X_22393_ _02800_ VPWR VGND _02897_ sg13g2_buf_1
X_22394_ _10631_ _02883_ VPWR VGND _02898_ sg13g2_nand2_1
X_22395_ _08694_ _02897_ _02898_ VPWR VGND _00419_ sg13g2_o21ai_1
X_22396_ _10633_ _02883_ VPWR VGND _02899_ sg13g2_nand2_1
X_22397_ _08715_ _02897_ _02899_ VPWR VGND _00420_ sg13g2_o21ai_1
X_22398_ _02775_ VPWR VGND _02900_ sg13g2_buf_1
X_22399_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[17]\ _02900_ VPWR VGND _02901_ sg13g2_nand2_1
X_22400_ _08714_ _02897_ _02901_ VPWR VGND _00421_ sg13g2_o21ai_1
X_22401_ _10285_ VPWR VGND _02902_ sg13g2_buf_1
X_22402_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ _02902_ VPWR VGND _00422_ sg13g2_mux2_1
X_22403_ _10723_ _10876_ _02902_ VPWR VGND _00423_ sg13g2_mux2_1
X_22404_ _10874_ _02900_ VPWR VGND _02903_ sg13g2_nand2_1
X_22405_ _10722_ _02897_ _02903_ VPWR VGND _00424_ sg13g2_o21ai_1
X_22406_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _02900_ VPWR VGND _02904_ sg13g2_nand2_1
X_22407_ _10721_ _02897_ _02904_ VPWR VGND _00425_ sg13g2_o21ai_1
X_22408_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _02900_ VPWR VGND _02905_ sg13g2_nand2_1
X_22409_ _08487_ _02897_ _02905_ VPWR VGND _00426_ sg13g2_o21ai_1
X_22410_ _10729_ _10871_ _02902_ VPWR VGND _00427_ sg13g2_mux2_1
X_22411_ _10736_ _10884_ _02902_ VPWR VGND _00428_ sg13g2_mux2_1
X_22412_ _10646_ _10885_ _02902_ VPWR VGND _00429_ sg13g2_mux2_1
X_22413_ _10647_ _10810_ _02902_ VPWR VGND _00430_ sg13g2_mux2_1
X_22414_ _10643_ _10807_ _02902_ VPWR VGND _00431_ sg13g2_mux2_1
X_22415_ _08759_ VPWR VGND _02906_ sg13g2_buf_1
X_22416_ _10642_ _02906_ VPWR VGND _02907_ sg13g2_nand2_1
X_22417_ _10816_ _02889_ _02907_ VPWR VGND _00432_ sg13g2_o21ai_1
X_22418_ _10652_ _10802_ _02902_ VPWR VGND _00433_ sg13g2_mux2_1
X_22419_ _10799_ _02900_ VPWR VGND _02908_ sg13g2_nand2_1
X_22420_ _10664_ _02897_ _02908_ VPWR VGND _00434_ sg13g2_o21ai_1
X_22421_ _10636_ _10800_ _02902_ VPWR VGND _00435_ sg13g2_mux2_1
X_22422_ _10635_ _02906_ VPWR VGND _02909_ sg13g2_nand2_1
X_22423_ _10833_ _02889_ _02909_ VPWR VGND _00436_ sg13g2_o21ai_1
X_22424_ _08483_ _02900_ VPWR VGND _02910_ sg13g2_nand2_1
X_22425_ _08884_ _02897_ _02910_ VPWR VGND _00437_ sg13g2_o21ai_1
X_22426_ _10676_ _10828_ _02902_ VPWR VGND _00438_ sg13g2_mux2_1
X_22427_ _10798_ _02900_ VPWR VGND _02911_ sg13g2_nand2_1
X_22428_ _10632_ _02897_ _02911_ VPWR VGND _00439_ sg13g2_o21ai_1
X_22429_ _10797_ _02900_ VPWR VGND _02912_ sg13g2_nand2_1
X_22430_ _10634_ _02897_ _02912_ VPWR VGND _00440_ sg13g2_o21ai_1
X_22431_ _02800_ VPWR VGND _02913_ sg13g2_buf_1
X_22432_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[17]\ _02900_ VPWR VGND _02914_ sg13g2_nand2_1
X_22433_ _10630_ _02913_ _02914_ VPWR VGND _00441_ sg13g2_o21ai_1
X_22434_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ _02896_ VPWR VGND _00442_ sg13g2_mux2_1
X_22435_ _11052_ _10876_ _02896_ VPWR VGND _00443_ sg13g2_mux2_1
X_22436_ _11050_ _10874_ _02896_ VPWR VGND _00444_ sg13g2_mux2_1
X_22437_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[60]\ _02900_ VPWR VGND _02915_ sg13g2_nand2_1
X_22438_ _10873_ _02913_ _02915_ VPWR VGND _00445_ sg13g2_o21ai_1
X_22439_ _10871_ _02906_ VPWR VGND _02916_ sg13g2_nand2_1
X_22440_ _11064_ _02889_ _02916_ VPWR VGND _00446_ sg13g2_o21ai_1
X_22441_ _10884_ _02906_ VPWR VGND _02917_ sg13g2_nand2_1
X_22442_ _11063_ _02889_ _02917_ VPWR VGND _00447_ sg13g2_o21ai_1
X_22443_ _02775_ VPWR VGND _02918_ sg13g2_buf_1
X_22444_ _08478_ _02918_ VPWR VGND _02919_ sg13g2_nand2_1
X_22445_ _09061_ _02913_ _02919_ VPWR VGND _00448_ sg13g2_o21ai_1
X_22446_ _10974_ _10885_ _02896_ VPWR VGND _00449_ sg13g2_mux2_1
X_22447_ _10975_ _10810_ _02896_ VPWR VGND _00450_ sg13g2_mux2_1
X_22448_ _10971_ _10807_ _02896_ VPWR VGND _00451_ sg13g2_mux2_1
X_22449_ _10970_ _02918_ VPWR VGND _02920_ sg13g2_nand2_1
X_22450_ _10816_ _02913_ _02920_ VPWR VGND _00452_ sg13g2_o21ai_1
X_22451_ _10981_ _10802_ _02896_ VPWR VGND _00453_ sg13g2_mux2_1
X_22452_ _10992_ _10799_ _02896_ VPWR VGND _00454_ sg13g2_mux2_1
X_22453_ _10991_ _10800_ _02896_ VPWR VGND _00455_ sg13g2_mux2_1
X_22454_ _10969_ _02918_ VPWR VGND _02921_ sg13g2_nand2_1
X_22455_ _10833_ _02913_ _02921_ VPWR VGND _00456_ sg13g2_o21ai_1
X_22456_ _10628_ VPWR VGND _02922_ sg13g2_buf_1
X_22457_ _10967_ _10828_ _02922_ VPWR VGND _00457_ sg13g2_mux2_1
X_22458_ _10798_ _02906_ VPWR VGND _02923_ sg13g2_nand2_1
X_22459_ _11114_ _02889_ _02923_ VPWR VGND _00458_ sg13g2_o21ai_1
X_22460_ _08427_ _02918_ VPWR VGND _02924_ sg13g2_nand2_1
X_22461_ _08907_ _02913_ _02924_ VPWR VGND _00459_ sg13g2_o21ai_1
X_22462_ _10963_ _10797_ _02922_ VPWR VGND _00460_ sg13g2_mux2_1
X_22463_ _11015_ _02918_ VPWR VGND _02925_ sg13g2_nand2_1
X_22464_ _10950_ _02913_ _02925_ VPWR VGND _00461_ sg13g2_o21ai_1
X_22465_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ _02922_ VPWR VGND _00462_ sg13g2_mux2_1
X_22466_ _11248_ _11052_ _02922_ VPWR VGND _00463_ sg13g2_mux2_1
X_22467_ _11246_ _11050_ _02922_ VPWR VGND _00464_ sg13g2_mux2_1
X_22468_ _11245_ _02918_ VPWR VGND _02926_ sg13g2_nand2_1
X_22469_ _11049_ _02913_ _02926_ VPWR VGND _00465_ sg13g2_o21ai_1
X_22470_ _11255_ _02918_ VPWR VGND _02927_ sg13g2_nand2_1
X_22471_ _11064_ _02913_ _02927_ VPWR VGND _00466_ sg13g2_o21ai_1
X_22472_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[81]\ _02918_ VPWR VGND _02928_ sg13g2_nand2_1
X_22473_ _11063_ _02913_ _02928_ VPWR VGND _00467_ sg13g2_o21ai_1
X_22474_ _11152_ _10974_ _02922_ VPWR VGND _00468_ sg13g2_mux2_1
X_22475_ _11153_ _10975_ _02922_ VPWR VGND _00469_ sg13g2_mux2_1
X_22476_ _08428_ _02918_ VPWR VGND _02929_ sg13g2_nand2_1
X_22477_ _12416_ _02774_ _02929_ VPWR VGND _00470_ sg13g2_o21ai_1
X_22478_ _11149_ _10971_ _02922_ VPWR VGND _00471_ sg13g2_mux2_1
X_22479_ _11148_ _02918_ VPWR VGND _02930_ sg13g2_nand2_1
X_22480_ _10986_ _02774_ _02930_ VPWR VGND _00472_ sg13g2_o21ai_1
X_22481_ _11159_ _10981_ _02922_ VPWR VGND _00473_ sg13g2_mux2_1
X_22482_ _10992_ _02906_ VPWR VGND _02931_ sg13g2_nand2_1
X_22483_ _11169_ _02889_ _02931_ VPWR VGND _00474_ sg13g2_o21ai_1
X_22484_ _11141_ _10991_ _02922_ VPWR VGND _00475_ sg13g2_mux2_1
X_22485_ _11140_ _10969_ _10619_ VPWR VGND _00476_ sg13g2_mux2_1
X_22486_ _11143_ _10967_ _10619_ VPWR VGND _00477_ sg13g2_mux2_1
X_22487_ _11180_ _11323_ VPWR VGND _02932_ sg13g2_nand2_1
X_22488_ _11114_ _02774_ _02932_ VPWR VGND _00478_ sg13g2_o21ai_1
X_22489_ _11138_ _10963_ _10619_ VPWR VGND _00479_ sg13g2_mux2_1
X_22490_ _11187_ _11015_ _10619_ VPWR VGND _00480_ sg13g2_mux2_1
X_22491_ _10586_ _08418_ _02776_ VPWR VGND _00481_ sg13g2_mux2_1
X_22492_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ _02776_ VPWR VGND _00482_ sg13g2_mux2_1
X_22493_ _11248_ _08890_ _02776_ VPWR VGND _00483_ sg13g2_mux2_1
X_22494_ _11246_ _02906_ VPWR VGND _02933_ sg13g2_nand2_1
X_22495_ _08887_ _02889_ _02933_ VPWR VGND _00484_ sg13g2_o21ai_1
X_22496_ _11245_ _02906_ VPWR VGND _02934_ sg13g2_nand2_1
X_22497_ _08886_ _02889_ _02934_ VPWR VGND _00485_ sg13g2_o21ai_1
X_22498_ _11255_ _02906_ VPWR VGND _02935_ sg13g2_nand2_1
X_22499_ _08881_ _09154_ _02935_ VPWR VGND _00486_ sg13g2_o21ai_1
X_22500_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _11323_ VPWR VGND _02936_ sg13g2_nand2_1
X_22501_ _11260_ _02774_ _02936_ VPWR VGND _00487_ sg13g2_o21ai_1
X_22502_ _11152_ _08771_ _02776_ VPWR VGND _00488_ sg13g2_mux2_1
X_22503_ _11153_ _08772_ _02776_ VPWR VGND _00489_ sg13g2_mux2_1
X_22504_ _11149_ _08769_ _02776_ VPWR VGND _00490_ sg13g2_mux2_1
X_22505_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[9]\ _11323_ VPWR VGND _02937_ sg13g2_nand2_1
X_22506_ _11211_ _02774_ _02937_ VPWR VGND _00491_ sg13g2_o21ai_1
X_22507_ _12404_ _02906_ VPWR VGND _02938_ sg13g2_nand2_1
X_22508_ _08444_ _09154_ _02938_ VPWR VGND _00492_ sg13g2_o21ai_1
X_22509_ _07679_ \atbs_core_0.dac_control_0.dac_init_value[1]\ VPWR VGND _02939_ sg13g2_nand2_1
X_22510_ _07679_ _11385_ _02939_ VPWR VGND _00545_ sg13g2_o21ai_1
X_22511_ _07679_ \atbs_core_0.dac_control_0.dac_init_value[2]\ VPWR VGND _02940_ sg13g2_nand2_1
X_22512_ _07679_ _11424_ _02940_ VPWR VGND _00546_ sg13g2_o21ai_1
X_22513_ _11382_ VPWR VGND _02941_ sg13g2_buf_1
X_22514_ _11416_ _02941_ VPWR VGND _02942_ sg13g2_nand2_1
X_22515_ _07678_ _07807_ _02942_ VPWR VGND _02943_ sg13g2_nor3_1
X_22516_ _07679_ \atbs_core_0.dac_control_0.dac_init_value[3]\ _02943_ VPWR VGND _00547_ sg13g2_a21o_1
X_22517_ _07678_ \atbs_core_0.dac_control_0.dac_init_value[4]\ VPWR VGND _02944_ sg13g2_nand2_1
X_22518_ _07679_ _11396_ _02944_ VPWR VGND _00548_ sg13g2_o21ai_1
X_22519_ _07678_ \atbs_core_0.dac_control_0.dac_init_value[5]\ VPWR VGND _02945_ sg13g2_nand2_1
X_22520_ _07679_ _11674_ _02945_ VPWR VGND _00549_ sg13g2_o21ai_1
X_22521_ \atbs_core_0.dac_control_0.dac_init_value[6]\ _07679_ VPWR VGND _00550_ sg13g2_nand2b_1
X_22522_ _07679_ \atbs_core_0.dac_control_0.dac_init_value[7]\ VPWR VGND _00551_ sg13g2_and2_1
X_22523_ \atbs_core_0.dac_control_1.dac_init_value[6]\ \atbs_core_0.dac_control_1.n1981_o\ VPWR VGND _00565_ sg13g2_nand2b_1
X_22524_ _07704_ _07705_ _07694_ _07703_ VPWR VGND 
+ _02946_
+ sg13g2_nor4_1
X_22525_ _02946_ _07903_ VPWR VGND _02947_ sg13g2_nor2b_1
X_22526_ _07909_ _07903_ _07655_ VPWR VGND _02948_ sg13g2_nor3_1
X_22527_ _07909_ _02947_ _02948_ VPWR VGND _02949_ sg13g2_a21oi_1
X_22528_ _07691_ _07693_ VPWR VGND _02950_ sg13g2_nand2_1
X_22529_ \atbs_core_0.main_counter_value[3]\ _02950_ _07707_ VPWR VGND _02951_ sg13g2_nor3_1
X_22530_ _07682_ _07905_ _02951_ VPWR VGND _02952_ sg13g2_nor3_1
X_22531_ _07709_ _07919_ _02952_ VPWR VGND _02953_ sg13g2_nor3_1
X_22532_ _07684_ _02949_ _02953_ VPWR VGND _02954_ sg13g2_o21ai_1
X_22533_ _07902_ _07914_ _07903_ VPWR VGND _02955_ sg13g2_a21oi_1
X_22534_ _07909_ _02955_ VPWR VGND _02956_ sg13g2_nor2_1
X_22535_ _07681_ _07686_ VPWR VGND _02957_ sg13g2_nand2_1
X_22536_ _12245_ _02956_ _02957_ VPWR VGND _02958_ sg13g2_nor3_1
X_22537_ _02954_ _02958_ VPWR VGND _00187_ sg13g2_nor2_1
X_22538_ _02734_ VPWR VGND _02959_ sg13g2_inv_1
X_22539_ _07675_ uart_rx_i _02959_ _07660_ VPWR VGND 
+ _00189_
+ sg13g2_a22oi_1
X_22540_ \atbs_core_0.memory2uart_0.n2605_q\ VPWR VGND _02960_ sg13g2_inv_1
X_22541_ _07649_ _07637_ VPWR VGND _02961_ sg13g2_and2_1
X_22542_ _07638_ _02960_ _02961_ _00062_ VPWR VGND 
+ _00190_
+ sg13g2_a22oi_1
X_22543_ _07996_ _07954_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1685_o\ sg13g2_nor2_1
X_22544_ _09534_ VPWR VGND _02962_ sg13g2_inv_1
X_22545_ _10288_ _10112_ VPWR VGND _02963_ sg13g2_nand2_1
X_22546_ _10450_ _10458_ VPWR VGND _02964_ sg13g2_nand2_1
X_22547_ _10289_ _10284_ VPWR VGND _02965_ sg13g2_nor2_1
X_22548_ _02964_ _02965_ VPWR VGND _02966_ sg13g2_nor2b_1
X_22549_ _00102_ VPWR VGND _02967_ sg13g2_buf_2
X_22550_ _10454_ _10450_ VPWR VGND _02968_ sg13g2_or2_1
X_22551_ _10622_ _02968_ _10458_ VPWR VGND _02969_ sg13g2_a21oi_1
X_22552_ _00103_ VPWR VGND _02970_ sg13g2_buf_2
X_22553_ _10454_ _10450_ _02970_ VPWR VGND _02971_ sg13g2_o21ai_1
X_22554_ _02971_ VPWR VGND _02972_ sg13g2_buf_1
X_22555_ _02972_ VPWR VGND _02973_ sg13g2_inv_1
X_22556_ _02967_ _02969_ _02973_ _02965_ VPWR VGND 
+ _02974_
+ sg13g2_or4_1
X_22557_ _02966_ _02974_ _10115_ VPWR VGND _02975_ sg13g2_nand3b_1
X_22558_ _10450_ VPWR VGND _02976_ sg13g2_inv_1
X_22559_ _10458_ _10621_ VPWR VGND _02977_ sg13g2_nor2b_1
X_22560_ _02977_ VPWR VGND _02978_ sg13g2_buf_2
X_22561_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2674_o[0]\ _02970_ VPWR VGND _02979_ sg13g2_and2_1
X_22562_ _02979_ VPWR VGND _02980_ sg13g2_buf_1
X_22563_ _02976_ _02978_ _02980_ VPWR VGND _02981_ sg13g2_a21oi_1
X_22564_ _10458_ _02970_ VPWR VGND _02982_ sg13g2_nor2b_1
X_22565_ _10455_ _02982_ _10284_ VPWR VGND _02983_ sg13g2_a21oi_1
X_22566_ _10455_ _02981_ _02983_ VPWR VGND _02984_ sg13g2_o21ai_1
X_22567_ _10450_ _10454_ VPWR VGND _02985_ sg13g2_nor2b_1
X_22568_ _02985_ VPWR VGND _02986_ sg13g2_buf_1
X_22569_ _02978_ _02986_ _02967_ VPWR VGND _02987_ sg13g2_a21oi_1
X_22570_ _10284_ _02987_ _10289_ VPWR VGND _02988_ sg13g2_a21oi_1
X_22571_ _10622_ _02968_ _10458_ VPWR VGND _02989_ sg13g2_a21o_1
X_22572_ _02989_ _02972_ _02987_ VPWR VGND _02990_ sg13g2_a21oi_1
X_22573_ _00101_ VPWR VGND _02991_ sg13g2_buf_1
X_22574_ _02984_ _02988_ _02990_ _10289_ _02991_ VPWR 
+ VGND
+ _02992_ sg13g2_a221oi_1
X_22575_ _02963_ _02975_ _02992_ VPWR VGND _02993_ sg13g2_a21o_1
X_22576_ _02993_ VPWR VGND _02994_ sg13g2_buf_1
X_22577_ _02967_ VPWR VGND _02995_ sg13g2_inv_1
X_22578_ _10455_ _10450_ _10621_ VPWR VGND _02996_ sg13g2_or3_1
X_22579_ _02970_ _10455_ VPWR VGND _02997_ sg13g2_nand2b_1
X_22580_ _10459_ _02996_ _02997_ VPWR VGND _02998_ sg13g2_nand3_1
X_22581_ _02995_ _02998_ VPWR VGND _02999_ sg13g2_nand2_1
X_22582_ _02970_ _02967_ _10459_ VPWR VGND _03000_ sg13g2_o21ai_1
X_22583_ _10450_ _03000_ VPWR VGND _03001_ sg13g2_nand2_1
X_22584_ _10289_ _02999_ _03001_ VPWR VGND _03002_ sg13g2_nand3_1
X_22585_ _03002_ VPWR VGND _03003_ sg13g2_buf_1
X_22586_ _10455_ VPWR VGND _03004_ sg13g2_inv_1
X_22587_ _02976_ _02978_ _02980_ VPWR VGND _03005_ sg13g2_a21o_1
X_22588_ _03004_ _10458_ VPWR VGND _03006_ sg13g2_nor2_1
X_22589_ _10284_ _02995_ VPWR VGND _03007_ sg13g2_nand2_1
X_22590_ _03004_ _03005_ _03006_ _02970_ _03007_ VPWR 
+ VGND
+ _03008_ sg13g2_a221oi_1
X_22591_ _10284_ _02969_ _02973_ VPWR VGND _03009_ sg13g2_nor3_1
X_22592_ _10289_ _03008_ _03009_ VPWR VGND _03010_ sg13g2_or3_1
X_22593_ _03010_ VPWR VGND _03011_ sg13g2_buf_2
X_22594_ _10288_ _10283_ VPWR VGND _03012_ sg13g2_nand2_1
X_22595_ _03003_ _03011_ _03012_ VPWR VGND _03013_ sg13g2_a21o_1
X_22596_ _03013_ VPWR VGND _03014_ sg13g2_buf_1
X_22597_ _02994_ _03014_ VPWR VGND _03015_ sg13g2_and2_1
X_22598_ _03015_ VPWR VGND _03016_ sg13g2_buf_1
X_22599_ _00104_ VPWR VGND _03017_ sg13g2_buf_1
X_22600_ _03017_ VPWR VGND _03018_ sg13g2_inv_1
X_22601_ _02978_ _02986_ VPWR VGND _03019_ sg13g2_nand2_1
X_22602_ _02995_ _03019_ _02989_ _02972_ _10453_ VPWR 
+ VGND
+ _03020_ sg13g2_a221oi_1
X_22603_ _02984_ _02988_ _03020_ VPWR VGND _03021_ sg13g2_a21o_1
X_22604_ _02991_ VPWR VGND _03022_ sg13g2_inv_1
X_22605_ _10289_ _10449_ _02978_ _02986_ VPWR VGND 
+ _03023_
+ sg13g2_nand4_1
X_22606_ _03023_ VPWR VGND _03024_ sg13g2_buf_1
X_22607_ _03022_ _03024_ VPWR VGND _03025_ sg13g2_and2_1
X_22608_ _10288_ _03025_ VPWR VGND _03026_ sg13g2_nor2_1
X_22609_ _03004_ _03005_ _03006_ _02970_ VPWR VGND 
+ _03027_
+ sg13g2_a22oi_1
X_22610_ _10289_ _02967_ VPWR VGND _03028_ sg13g2_nand2_1
X_22611_ _10284_ _02967_ VPWR VGND _03029_ sg13g2_nand2_1
X_22612_ _10449_ _02978_ _02986_ VPWR VGND _03030_ sg13g2_nand3_1
X_22613_ _03029_ _03030_ _10289_ VPWR VGND _03031_ sg13g2_a21o_1
X_22614_ _03027_ _03028_ _03031_ VPWR VGND _03032_ sg13g2_o21ai_1
X_22615_ _03032_ VPWR VGND _03033_ sg13g2_buf_1
X_22616_ _10115_ _10112_ VPWR VGND _03034_ sg13g2_nor2_1
X_22617_ _03025_ _02963_ VPWR VGND _03035_ sg13g2_nor2_1
X_22618_ _03021_ _03026_ _03033_ _03034_ _03035_ VPWR 
+ VGND
+ _03036_ sg13g2_a221oi_1
X_22619_ _03036_ VPWR VGND _03037_ sg13g2_buf_2
X_22620_ _03018_ _03037_ VPWR VGND _03038_ sg13g2_nand2_1
X_22621_ _03016_ _03038_ VPWR VGND _03039_ sg13g2_nand2b_1
X_22622_ _09913_ _09712_ VPWR VGND _03040_ sg13g2_nor2_1
X_22623_ _03029_ _03030_ VPWR VGND _03041_ sg13g2_nand2_1
X_22624_ _10453_ _02995_ VPWR VGND _03042_ sg13g2_nor2_1
X_22625_ _10455_ _02982_ VPWR VGND _03043_ sg13g2_nand2_1
X_22626_ _10455_ _02981_ _03043_ VPWR VGND _03044_ sg13g2_o21ai_1
X_22627_ _10453_ _03041_ _03042_ _03044_ VPWR VGND 
+ _03045_
+ sg13g2_a22oi_1
X_22628_ _03022_ _03045_ _02963_ VPWR VGND _03046_ sg13g2_a21oi_1
X_22629_ _02984_ _02988_ _03020_ VPWR VGND _03047_ sg13g2_a21oi_1
X_22630_ _03047_ _03012_ VPWR VGND _03048_ sg13g2_nor2_1
X_22631_ _03022_ _03045_ _03003_ _03011_ _10288_ VPWR 
+ VGND
+ _03049_ sg13g2_a221oi_1
X_22632_ _03046_ _03048_ _03049_ VPWR VGND _03050_ sg13g2_or3_1
X_22633_ _03050_ VPWR VGND _03051_ sg13g2_buf_1
X_22634_ _03051_ VPWR VGND _03052_ sg13g2_inv_1
X_22635_ _09913_ VPWR VGND _03053_ sg13g2_inv_1
X_22636_ _03053_ _09712_ VPWR VGND _03054_ sg13g2_nand2_1
X_22637_ _03038_ _03054_ VPWR VGND _03055_ sg13g2_nor2_1
X_22638_ _09914_ _03039_ _03040_ _03052_ _03055_ VPWR 
+ VGND
+ _03056_ sg13g2_a221oi_1
X_22639_ _03056_ VPWR VGND _03057_ sg13g2_buf_1
X_22640_ _10288_ _03022_ VPWR VGND _03058_ sg13g2_nor2_1
X_22641_ _10112_ _02991_ VPWR VGND _03059_ sg13g2_nand2_1
X_22642_ _10112_ _03024_ _03059_ VPWR VGND _03060_ sg13g2_o21ai_1
X_22643_ _10288_ _03060_ VPWR VGND _03061_ sg13g2_and2_1
X_22644_ _03033_ _03058_ _03061_ VPWR VGND _03062_ sg13g2_a21o_1
X_22645_ _09712_ _03018_ VPWR VGND _03063_ sg13g2_nand2_1
X_22646_ _09712_ _03062_ _03063_ VPWR VGND _03064_ sg13g2_o21ai_1
X_22647_ _03037_ _03017_ _09914_ VPWR VGND _03065_ sg13g2_nand3b_1
X_22648_ _09914_ _03064_ _03065_ VPWR VGND _03066_ sg13g2_o21ai_1
X_22649_ _00105_ VPWR VGND _03067_ sg13g2_buf_1
X_22650_ _03067_ VPWR VGND _03068_ sg13g2_inv_1
X_22651_ _03066_ _03068_ VPWR VGND _03069_ sg13g2_nand2b_1
X_22652_ _09706_ _03057_ _03069_ VPWR VGND _03070_ sg13g2_and3_1
X_22653_ _09706_ _09537_ VPWR VGND _03071_ sg13g2_nand2b_1
X_22654_ _03071_ _03069_ VPWR VGND _03072_ sg13g2_nor2b_1
X_22655_ _09712_ VPWR VGND _03073_ sg13g2_inv_1
X_22656_ _03033_ _03058_ VPWR VGND _03074_ sg13g2_nand2_1
X_22657_ _03061_ _03063_ VPWR VGND _03075_ sg13g2_nor2_1
X_22658_ _03073_ _03037_ _03074_ _03075_ VPWR VGND 
+ _03076_
+ sg13g2_a22oi_1
X_22659_ _10288_ _03060_ _03058_ _03033_ _03017_ VPWR 
+ VGND
+ _03077_ sg13g2_a221oi_1
X_22660_ _03053_ _03077_ VPWR VGND _03078_ sg13g2_nor2_1
X_22661_ _03053_ _03076_ _03051_ _03078_ VPWR VGND 
+ _03079_
+ sg13g2_a22oi_1
X_22662_ _03079_ VPWR VGND _03080_ sg13g2_buf_1
X_22663_ _09706_ _09537_ VPWR VGND _03081_ sg13g2_nor2_1
X_22664_ _03081_ VPWR VGND _03082_ sg13g2_buf_1
X_22665_ _03080_ _03082_ VPWR VGND _03083_ sg13g2_nor2b_1
X_22666_ _03070_ _03072_ _03083_ VPWR VGND _03084_ sg13g2_nor3_1
X_22667_ _00106_ VPWR VGND _03085_ sg13g2_buf_1
X_22668_ _03085_ VPWR VGND _03086_ sg13g2_inv_1
X_22669_ _09537_ _03068_ VPWR VGND _03087_ sg13g2_nand2_1
X_22670_ _09537_ _03066_ _03087_ VPWR VGND _03088_ sg13g2_o21ai_1
X_22671_ _03080_ _03067_ VPWR VGND _03089_ sg13g2_nand2b_1
X_22672_ _03088_ _03089_ _09706_ VPWR VGND _03090_ sg13g2_mux2_1
X_22673_ _03090_ VPWR VGND _03091_ sg13g2_buf_1
X_22674_ _09533_ _09342_ VPWR VGND _03092_ sg13g2_nor2_1
X_22675_ _03086_ _03091_ _03092_ VPWR VGND _03093_ sg13g2_a21oi_1
X_22676_ _03093_ VPWR VGND _03094_ sg13g2_inv_1
X_22677_ _09342_ _03084_ _03094_ VPWR VGND _03095_ sg13g2_o21ai_1
X_22678_ _03063_ _03046_ _03048_ _03049_ VPWR VGND 
+ _03096_
+ sg13g2_or4_1
X_22679_ _03073_ _02994_ _03014_ VPWR VGND _03097_ sg13g2_nand3_1
X_22680_ _03053_ _03096_ _03097_ VPWR VGND _03098_ sg13g2_nand3_1
X_22681_ _03098_ VPWR VGND _03099_ sg13g2_buf_1
X_22682_ _03017_ _03046_ _03048_ _03049_ VPWR VGND 
+ _03100_
+ sg13g2_or4_1
X_22683_ _02995_ _02998_ _03000_ _10450_ _10453_ VPWR 
+ VGND
+ _03101_ sg13g2_a221oi_1
X_22684_ _02991_ _03101_ VPWR VGND _03102_ sg13g2_nor2_1
X_22685_ _02967_ _02964_ _02965_ VPWR VGND _03103_ sg13g2_or3_1
X_22686_ _03103_ VPWR VGND _03104_ sg13g2_buf_1
X_22687_ _10115_ _03104_ VPWR VGND _03105_ sg13g2_nand2_1
X_22688_ _03011_ _03102_ _03105_ VPWR VGND _03106_ sg13g2_a21oi_1
X_22689_ _02966_ _02974_ VPWR VGND _03107_ sg13g2_nand2b_1
X_22690_ _03107_ VPWR VGND _03108_ sg13g2_buf_1
X_22691_ _10283_ _02991_ _03101_ VPWR VGND _03109_ sg13g2_nor3_1
X_22692_ _10283_ _03108_ _03109_ _03011_ _10115_ VPWR 
+ VGND
+ _03110_ sg13g2_a221oi_1
X_22693_ _03106_ _03110_ VPWR VGND _03111_ sg13g2_or2_1
X_22694_ _03111_ VPWR VGND _03112_ sg13g2_buf_1
X_22695_ _09914_ _03100_ _03112_ VPWR VGND _03113_ sg13g2_nand3_1
X_22696_ _03113_ VPWR VGND _03114_ sg13g2_buf_1
X_22697_ _03068_ _03080_ _03099_ _03114_ VPWR VGND 
+ _03115_
+ sg13g2_a22oi_1
X_22698_ _03068_ _03080_ _03071_ VPWR VGND _03116_ sg13g2_a21oi_1
X_22699_ _03057_ _03082_ _03115_ _09706_ _03116_ VPWR 
+ VGND
+ _03117_ sg13g2_a221oi_1
X_22700_ _03117_ VPWR VGND _03118_ sg13g2_buf_1
X_22701_ _03118_ VPWR VGND _03119_ sg13g2_inv_1
X_22702_ _02962_ _03095_ _03119_ _03093_ VPWR VGND 
+ _03120_
+ sg13g2_a22oi_1
X_22703_ _09340_ _03120_ VPWR VGND _03121_ sg13g2_nor2_1
X_22704_ _03086_ _03084_ VPWR VGND _03122_ sg13g2_nor2_1
X_22705_ _03085_ _09342_ VPWR VGND _03123_ sg13g2_nor2b_1
X_22706_ _09342_ _03091_ VPWR VGND _03124_ sg13g2_nor2b_1
X_22707_ _09534_ _03123_ _03124_ VPWR VGND _03125_ sg13g2_nor3_1
X_22708_ _09534_ _03122_ _03125_ VPWR VGND _03126_ sg13g2_a21oi_1
X_22709_ _09339_ _03126_ VPWR VGND _03127_ sg13g2_nor2_1
X_22710_ _03121_ _03127_ _09337_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[48]\ sg13g2_o21ai_1
X_22711_ _09339_ _09336_ VPWR VGND _03128_ sg13g2_nor2_1
X_22712_ _09336_ _03126_ _03128_ _03120_ VPWR VGND 
+ _03129_
+ sg13g2_a22oi_1
X_22713_ _09537_ _03099_ _03114_ VPWR VGND _03130_ sg13g2_nand3b_1
X_22714_ _03018_ _03037_ _02994_ _03014_ VPWR VGND 
+ _03131_
+ sg13g2_a22oi_1
X_22715_ _03018_ _03037_ _03054_ VPWR VGND _03132_ sg13g2_a21oi_1
X_22716_ _09914_ _03131_ _03132_ VPWR VGND _03133_ sg13g2_a21oi_1
X_22717_ _03051_ _03040_ _03087_ VPWR VGND _03134_ sg13g2_a21oi_1
X_22718_ _03133_ _03134_ _09706_ VPWR VGND _03135_ sg13g2_a21oi_1
X_22719_ _02967_ _02964_ _02965_ VPWR VGND _03136_ sg13g2_nor3_1
X_22720_ _02991_ _03034_ VPWR VGND _03137_ sg13g2_nor2_1
X_22721_ _03034_ _03136_ _03137_ _03108_ VPWR VGND 
+ _03138_
+ sg13g2_a22oi_1
X_22722_ _09913_ _03138_ VPWR VGND _03139_ sg13g2_nand2_1
X_22723_ _03018_ _03016_ _03054_ _03139_ VPWR VGND 
+ _03140_
+ sg13g2_a22oi_1
X_22724_ _03040_ _03112_ VPWR VGND _03141_ sg13g2_and2_1
X_22725_ _03140_ _03141_ VPWR VGND _03142_ sg13g2_or2_1
X_22726_ _03142_ VPWR VGND _03143_ sg13g2_buf_1
X_22727_ _09914_ _09712_ _03067_ VPWR VGND _03144_ sg13g2_nor3_1
X_22728_ _03053_ _03067_ VPWR VGND _03145_ sg13g2_nor2_1
X_22729_ _03053_ _09712_ _03068_ VPWR VGND _03146_ sg13g2_nand3_1
X_22730_ _03038_ _03146_ _09706_ VPWR VGND _03147_ sg13g2_o21ai_1
X_22731_ _03052_ _03144_ _03145_ _03039_ _03147_ VPWR 
+ VGND
+ _03148_ sg13g2_a221oi_1
X_22732_ _03130_ _03135_ _03143_ _03148_ VPWR VGND 
+ _03149_
+ sg13g2_a22oi_1
X_22733_ _03086_ _03084_ _03149_ _09534_ _03092_ VPWR 
+ VGND
+ _03150_ sg13g2_a221oi_1
X_22734_ _03092_ _03119_ _03150_ VPWR VGND _03151_ sg13g2_a21oi_1
X_22735_ _09339_ _03151_ VPWR VGND _03152_ sg13g2_nand2_1
X_22736_ _03129_ _03152_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[49]\ sg13g2_nand2_1
X_22737_ _09336_ _03120_ _03128_ _03151_ VPWR VGND 
+ _03153_
+ sg13g2_a22oi_1
X_22738_ _03086_ _03118_ VPWR VGND _03154_ sg13g2_nand2_1
X_22739_ _03012_ _03104_ VPWR VGND _03155_ sg13g2_nor2_1
X_22740_ _03108_ _03137_ _03155_ VPWR VGND _03156_ sg13g2_a21o_1
X_22741_ _03017_ _03040_ VPWR VGND _03157_ sg13g2_nor2_1
X_22742_ _03106_ _03110_ VPWR VGND _03158_ sg13g2_nor2_1
X_22743_ _03040_ _03156_ _03157_ _03158_ VPWR VGND 
+ _03159_
+ sg13g2_a22oi_1
X_22744_ _09706_ _03159_ VPWR VGND _03160_ sg13g2_nand2_1
X_22745_ _03068_ _03099_ _03114_ VPWR VGND _03161_ sg13g2_and3_1
X_22746_ _03071_ _03160_ _03161_ VPWR VGND _03162_ sg13g2_a21oi_1
X_22747_ _03082_ _03143_ _03162_ VPWR VGND _03163_ sg13g2_a21o_1
X_22748_ _03163_ VPWR VGND _03164_ sg13g2_buf_1
X_22749_ _09534_ _03154_ _03164_ VPWR VGND _03165_ sg13g2_nand3_1
X_22750_ _09533_ _09342_ VPWR VGND _03166_ sg13g2_nor2b_1
X_22751_ _09533_ _09342_ VPWR VGND _03167_ sg13g2_or2_1
X_22752_ _03167_ VPWR VGND _03168_ sg13g2_buf_1
X_22753_ _03168_ _03149_ VPWR VGND _03169_ sg13g2_nor2_1
X_22754_ _03154_ _03166_ _03169_ VPWR VGND _03170_ sg13g2_a21oi_1
X_22755_ _03165_ _03170_ VPWR VGND _03171_ sg13g2_and2_1
X_22756_ _03171_ VPWR VGND _03172_ sg13g2_buf_1
X_22757_ _09339_ _03172_ VPWR VGND _03173_ sg13g2_nand2_1
X_22758_ _03153_ _03173_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[50]\ sg13g2_nand2_1
X_22759_ _03082_ _03143_ _03162_ VPWR VGND _03174_ sg13g2_a21oi_1
X_22760_ _03130_ _03135_ _03143_ _03148_ _03085_ VPWR 
+ VGND
+ _03175_ sg13g2_a221oi_1
X_22761_ _03067_ _03140_ _03141_ VPWR VGND _03176_ sg13g2_nor3_1
X_22762_ _03082_ _03159_ VPWR VGND _03177_ sg13g2_nand2_1
X_22763_ _03082_ _03176_ _03177_ VPWR VGND _03178_ sg13g2_o21ai_1
X_22764_ _03175_ _03178_ VPWR VGND _03179_ sg13g2_nor2b_1
X_22765_ _03175_ _03166_ VPWR VGND _03180_ sg13g2_nor2b_1
X_22766_ _09534_ _03179_ _03180_ VPWR VGND _03181_ sg13g2_a21oi_1
X_22767_ _03168_ _03174_ _03181_ VPWR VGND _03182_ sg13g2_o21ai_1
X_22768_ _03182_ VPWR VGND _03183_ sg13g2_buf_1
X_22769_ _09336_ _03151_ _03172_ _03128_ VPWR VGND 
+ _03184_
+ sg13g2_a22oi_1
X_22770_ _09340_ _03183_ _03184_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[51]\ sg13g2_o21ai_1
X_22771_ _03128_ VPWR VGND _03185_ sg13g2_inv_1
X_22772_ _03168_ _03178_ VPWR VGND _03186_ sg13g2_nor2_1
X_22773_ _09342_ _03174_ _03186_ VPWR VGND _03187_ sg13g2_a21o_1
X_22774_ _03187_ VPWR VGND _03188_ sg13g2_buf_1
X_22775_ _09336_ _03172_ _03188_ _09339_ VPWR VGND 
+ _03189_
+ sg13g2_a22oi_1
X_22776_ _03185_ _03183_ _03189_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[52]\ sg13g2_o21ai_1
X_22777_ _03128_ _03188_ VPWR VGND _03190_ sg13g2_nand2_1
X_22778_ _09337_ _03183_ _03190_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[53]\ sg13g2_o21ai_1
X_22779_ _03092_ _03164_ _03179_ _09534_ _03180_ VPWR 
+ VGND
+ _03191_ sg13g2_a221oi_1
X_22780_ _09150_ _08979_ _00044_ VPWR VGND _03192_ sg13g2_nor3_1
X_22781_ _08980_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _09150_ VPWR VGND 
+ _03193_
+ sg13g2_a22oi_1
X_22782_ _03192_ _03193_ VPWR VGND _03194_ sg13g2_nand2b_1
X_22783_ _08972_ VPWR VGND _03195_ sg13g2_buf_2
X_22784_ _03195_ _08827_ VPWR VGND _03196_ sg13g2_nor2_1
X_22785_ _09150_ _08979_ VPWR VGND _03197_ sg13g2_or2_1
X_22786_ _03197_ VPWR VGND _03198_ sg13g2_buf_1
X_22787_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ VPWR VGND _03199_ sg13g2_buf_1
X_22788_ _08980_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ _03199_ _09150_ VPWR VGND 
+ _03200_
+ sg13g2_a22oi_1
X_22789_ _00046_ _03198_ _03200_ VPWR VGND _03201_ sg13g2_o21ai_1
X_22790_ _03201_ VPWR VGND _03202_ sg13g2_buf_2
X_22791_ _08980_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _09150_ VPWR VGND 
+ _03203_
+ sg13g2_a22oi_1
X_22792_ _09150_ _08980_ _00048_ VPWR VGND _03204_ sg13g2_or3_1
X_22793_ _03204_ VPWR VGND _03205_ sg13g2_buf_1
X_22794_ _03203_ _03205_ _08973_ VPWR VGND _03206_ sg13g2_a21oi_1
X_22795_ _08827_ _03194_ _03196_ _03202_ _03206_ VPWR 
+ VGND
+ _03207_ sg13g2_a221oi_1
X_22796_ _03207_ VPWR VGND _03208_ sg13g2_buf_1
X_22797_ _11135_ _03208_ VPWR VGND _03209_ sg13g2_nor2_1
X_22798_ _08974_ VPWR VGND _03210_ sg13g2_inv_1
X_22799_ _03210_ _11135_ VPWR VGND _03211_ sg13g2_nand2_1
X_22800_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ VPWR VGND _03212_ sg13g2_inv_1
X_22801_ _08980_ _03199_ VPWR VGND _03213_ sg13g2_nand2_1
X_22802_ _03212_ _03198_ _03213_ VPWR VGND _03214_ sg13g2_o21ai_1
X_22803_ _03195_ _08826_ VPWR VGND _03215_ sg13g2_or2_1
X_22804_ _03203_ _03205_ _03215_ VPWR VGND _03216_ sg13g2_a21oi_1
X_22805_ _08827_ _03202_ _03214_ _03195_ _03216_ VPWR 
+ VGND
+ _03217_ sg13g2_a221oi_1
X_22806_ _03217_ VPWR VGND _03218_ sg13g2_buf_1
X_22807_ _03211_ _03218_ VPWR VGND _03219_ sg13g2_nor2_1
X_22808_ _03203_ _03205_ VPWR VGND _03220_ sg13g2_nand2_1
X_22809_ _08827_ _03220_ _03214_ _03196_ VPWR VGND 
+ _03221_
+ sg13g2_a22oi_1
X_22810_ _03210_ _03221_ VPWR VGND _03222_ sg13g2_nor2_1
X_22811_ _03209_ _03219_ _03222_ VPWR VGND _03223_ sg13g2_or3_1
X_22812_ _03223_ VPWR VGND _03224_ sg13g2_buf_1
X_22813_ _03218_ _08756_ VPWR VGND _03225_ sg13g2_nand2b_1
X_22814_ _03211_ _03221_ VPWR VGND _03226_ sg13g2_or2_1
X_22815_ _11132_ _11123_ VPWR VGND _03227_ sg13g2_or2_1
X_22816_ _03227_ VPWR VGND _03228_ sg13g2_buf_1
X_22817_ _03225_ _03226_ _03228_ VPWR VGND _03229_ sg13g2_a21oi_1
X_22818_ _11123_ _03224_ _03229_ VPWR VGND _03230_ sg13g2_a21o_1
X_22819_ _03230_ VPWR VGND _03231_ sg13g2_buf_1
X_22820_ _10960_ _10957_ VPWR VGND _03232_ sg13g2_nor2_1
X_22821_ _10957_ VPWR VGND _03233_ sg13g2_inv_1
X_22822_ _03208_ _03211_ VPWR VGND _03234_ sg13g2_nor2_1
X_22823_ _03210_ _03218_ VPWR VGND _03235_ sg13g2_nor2_1
X_22824_ _03192_ _03193_ VPWR VGND _03236_ sg13g2_nor2b_1
X_22825_ _08979_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ _09149_ VPWR VGND 
+ _03237_
+ sg13g2_a22oi_1
X_22826_ _03237_ VPWR VGND _03238_ sg13g2_buf_1
X_22827_ _09149_ _08979_ _00042_ VPWR VGND _03239_ sg13g2_or3_1
X_22828_ _03239_ VPWR VGND _03240_ sg13g2_buf_1
X_22829_ _00041_ VPWR VGND _03241_ sg13g2_buf_1
X_22830_ _03238_ _03240_ _03241_ VPWR VGND _03242_ sg13g2_a21o_1
X_22831_ _03242_ VPWR VGND _03243_ sg13g2_buf_1
X_22832_ _03236_ _03243_ _08827_ VPWR VGND _03244_ sg13g2_mux2_1
X_22833_ _08973_ _03202_ VPWR VGND _03245_ sg13g2_nor2_1
X_22834_ _08973_ _03244_ _03245_ _03243_ _11135_ VPWR 
+ VGND
+ _03246_ sg13g2_a221oi_1
X_22835_ _03234_ _03235_ _03246_ VPWR VGND _03247_ sg13g2_or3_1
X_22836_ _03247_ VPWR VGND _03248_ sg13g2_buf_1
X_22837_ _11132_ _11123_ VPWR VGND _03249_ sg13g2_nor2_1
X_22838_ _03225_ _03226_ _11316_ VPWR VGND _03250_ sg13g2_a21oi_1
X_22839_ _11123_ _03248_ _03224_ _03249_ _03250_ VPWR 
+ VGND
+ _03251_ sg13g2_a221oi_1
X_22840_ _03251_ VPWR VGND _03252_ sg13g2_buf_1
X_22841_ _03233_ _03252_ VPWR VGND _03253_ sg13g2_nor2_1
X_22842_ _03231_ _03232_ _03253_ VPWR VGND _03254_ sg13g2_a21o_1
X_22843_ _03254_ VPWR VGND _03255_ sg13g2_buf_1
X_22844_ _03249_ _03248_ _03224_ _11132_ VPWR VGND 
+ _03256_
+ sg13g2_a22oi_1
X_22845_ _03241_ VPWR VGND _03257_ sg13g2_inv_1
X_22846_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ _09150_ VPWR VGND _03258_ sg13g2_nand2b_1
X_22847_ _09149_ _00040_ VPWR VGND _03259_ sg13g2_nand2b_1
X_22848_ _03258_ _03259_ _08979_ VPWR VGND _03260_ sg13g2_a21o_1
X_22849_ _03260_ VPWR VGND _03261_ sg13g2_buf_1
X_22850_ _08827_ _03257_ _03261_ VPWR VGND _03262_ sg13g2_nand3_1
X_22851_ _03262_ VPWR VGND _03263_ sg13g2_buf_1
X_22852_ _03238_ _03240_ _08827_ VPWR VGND _03264_ sg13g2_a21oi_1
X_22853_ _03195_ _03264_ VPWR VGND _03265_ sg13g2_nor2_1
X_22854_ _03257_ _03261_ _03194_ VPWR VGND _03266_ sg13g2_a21oi_1
X_22855_ _00043_ VPWR VGND _03267_ sg13g2_buf_1
X_22856_ _03267_ _08756_ VPWR VGND _03268_ sg13g2_nand2b_1
X_22857_ _03263_ _03265_ _03266_ _03195_ _03268_ VPWR 
+ VGND
+ _03269_ sg13g2_a221oi_1
X_22858_ _03267_ _08974_ VPWR VGND _03270_ sg13g2_nand2b_1
X_22859_ _03263_ _03265_ _03266_ _03195_ _03270_ VPWR 
+ VGND
+ _03271_ sg13g2_a221oi_1
X_22860_ _08973_ _03244_ _03245_ _03243_ _03211_ VPWR 
+ VGND
+ _03272_ sg13g2_a221oi_1
X_22861_ _03210_ _03208_ VPWR VGND _03273_ sg13g2_nor2_1
X_22862_ _03269_ _03271_ _03272_ _03273_ VPWR VGND 
+ _03274_
+ sg13g2_or4_1
X_22863_ _03274_ VPWR VGND _03275_ sg13g2_buf_1
X_22864_ _11123_ _03275_ VPWR VGND _03276_ sg13g2_nand2_1
X_22865_ _10960_ VPWR VGND _03277_ sg13g2_inv_1
X_22866_ _03277_ _03233_ VPWR VGND _03278_ sg13g2_nand2_1
X_22867_ _03256_ _03276_ _03278_ VPWR VGND _03279_ sg13g2_a21o_1
X_22868_ _03252_ _10960_ VPWR VGND _03280_ sg13g2_nand2b_1
X_22869_ _03192_ _03193_ _03195_ VPWR VGND _03281_ sg13g2_nand3b_1
X_22870_ _03257_ _03261_ _03281_ VPWR VGND _03282_ sg13g2_a21oi_1
X_22871_ _03263_ _03265_ _03282_ VPWR VGND _03283_ sg13g2_a21oi_1
X_22872_ _03195_ _08826_ _08980_ VPWR VGND _03284_ sg13g2_or3_1
X_22873_ _03258_ _03259_ _03284_ VPWR VGND _03285_ sg13g2_a21oi_1
X_22874_ _08973_ _08827_ _03241_ VPWR VGND _03286_ sg13g2_and3_1
X_22875_ _03286_ VPWR VGND _03287_ sg13g2_buf_1
X_22876_ _03195_ _03241_ _03238_ _03240_ VPWR VGND 
+ _03288_
+ sg13g2_and4_1
X_22877_ _03288_ VPWR VGND _03289_ sg13g2_buf_1
X_22878_ _03267_ _03285_ _03287_ _03289_ VPWR VGND 
+ _03290_
+ sg13g2_or4_1
X_22879_ _11135_ _03290_ _03210_ VPWR VGND _03291_ sg13g2_o21ai_1
X_22880_ _11135_ _03283_ _03291_ VPWR VGND _03292_ sg13g2_a21o_1
X_22881_ _03292_ VPWR VGND _03293_ sg13g2_buf_1
X_22882_ _03202_ _03243_ VPWR VGND _03294_ sg13g2_nor2b_1
X_22883_ _03244_ _03294_ _03195_ VPWR VGND _03295_ sg13g2_mux2_1
X_22884_ _03295_ VPWR VGND _03296_ sg13g2_buf_1
X_22885_ _08974_ _03290_ VPWR VGND _03297_ sg13g2_and2_1
X_22886_ _03296_ _03297_ _00045_ VPWR VGND _03298_ sg13g2_a21oi_1
X_22887_ _11316_ _11123_ VPWR VGND _03299_ sg13g2_nand2_1
X_22888_ _11316_ _03234_ _03235_ _03246_ VPWR VGND 
+ _03300_
+ sg13g2_or4_1
X_22889_ _03293_ _03298_ _03299_ _03300_ VPWR VGND 
+ _03301_
+ sg13g2_a22oi_1
X_22890_ _03228_ _03275_ VPWR VGND _03302_ sg13g2_nor2_1
X_22891_ _03233_ _03301_ _03302_ VPWR VGND _03303_ sg13g2_or3_1
X_22892_ _03279_ _03280_ _03303_ VPWR VGND _03304_ sg13g2_nand3_1
X_22893_ _03304_ VPWR VGND _03305_ sg13g2_buf_1
X_22894_ _10794_ _03255_ _03305_ _10624_ VPWR VGND 
+ _03306_
+ sg13g2_a22oi_1
X_22895_ _03256_ _03276_ _03233_ VPWR VGND _03307_ sg13g2_a21o_1
X_22896_ _10960_ _03231_ VPWR VGND _03308_ sg13g2_nand2_1
X_22897_ _03252_ _03232_ VPWR VGND _03309_ sg13g2_nand2b_1
X_22898_ _03307_ _03308_ _03309_ VPWR VGND _03310_ sg13g2_nand3_1
X_22899_ _03310_ VPWR VGND _03311_ sg13g2_buf_1
X_22900_ _10794_ _10624_ VPWR VGND _03312_ sg13g2_nor2_1
X_22901_ _03312_ VPWR VGND _03313_ sg13g2_buf_1
X_22902_ _09709_ _03313_ _03255_ VPWR VGND _03314_ sg13g2_and3_1
X_22903_ _02976_ _10459_ VPWR VGND _03315_ sg13g2_nor2_1
X_22904_ _03199_ _03315_ _03220_ VPWR VGND _03316_ sg13g2_nor3_1
X_22905_ _03218_ _03316_ VPWR VGND _03317_ sg13g2_nand2_1
X_22906_ _03108_ _03224_ _03317_ VPWR VGND _03318_ sg13g2_nor3_1
X_22907_ _03112_ _03143_ _03252_ _03318_ VPWR VGND 
+ _03319_
+ sg13g2_nand4_1
X_22908_ _03311_ _03314_ _03319_ VPWR VGND _03320_ sg13g2_nor3_1
X_22909_ _03164_ _03306_ _03320_ VPWR VGND _03321_ sg13g2_and3_1
X_22910_ _03256_ _03276_ VPWR VGND _03322_ sg13g2_nand2_1
X_22911_ _03263_ _03265_ _03282_ VPWR VGND _03323_ sg13g2_a21o_1
X_22912_ _03323_ VPWR VGND _03324_ sg13g2_buf_1
X_22913_ _08756_ _03208_ _08974_ VPWR VGND _03325_ sg13g2_mux2_1
X_22914_ _03267_ _03324_ _03325_ VPWR VGND _03326_ sg13g2_o21ai_1
X_22915_ _08974_ _08756_ VPWR VGND _03327_ sg13g2_nor2_1
X_22916_ _03327_ _03296_ _11316_ VPWR VGND _03328_ sg13g2_a21oi_1
X_22917_ _08974_ _03267_ VPWR VGND _03329_ sg13g2_and2_1
X_22918_ _03285_ _03287_ _03289_ VPWR VGND _03330_ sg13g2_nor3_1
X_22919_ _03210_ _03268_ VPWR VGND _03331_ sg13g2_nand2_1
X_22920_ _11135_ _03330_ _03331_ VPWR VGND _03332_ sg13g2_a21oi_1
X_22921_ _03324_ _03329_ _03332_ VPWR VGND _03333_ sg13g2_a21oi_1
X_22922_ _00045_ VPWR VGND _03334_ sg13g2_inv_1
X_22923_ _03326_ _03328_ _03333_ _03334_ _03249_ VPWR 
+ VGND
+ _03335_ sg13g2_a221oi_1
X_22924_ _03335_ VPWR VGND _03336_ sg13g2_buf_1
X_22925_ _03296_ _03297_ VPWR VGND _03337_ sg13g2_nand2_1
X_22926_ _03293_ _03337_ _03228_ VPWR VGND _03338_ sg13g2_a21oi_1
X_22927_ _00047_ _03336_ _03338_ VPWR VGND _03339_ sg13g2_nor3_1
X_22928_ _03277_ _03322_ _03339_ VPWR VGND _03340_ sg13g2_or3_1
X_22929_ _03340_ VPWR VGND _03341_ sg13g2_buf_1
X_22930_ _10957_ _03301_ _03302_ VPWR VGND _03342_ sg13g2_nor3_1
X_22931_ _03233_ _00047_ _03336_ _03338_ VPWR VGND 
+ _03343_
+ sg13g2_nor4_1
X_22932_ _10960_ _03342_ _03343_ VPWR VGND _03344_ sg13g2_or3_1
X_22933_ _03344_ VPWR VGND _03345_ sg13g2_buf_1
X_22934_ _10624_ _03341_ _03345_ VPWR VGND _03346_ sg13g2_nand3_1
X_22935_ _10794_ _03311_ _03313_ _03305_ VPWR VGND 
+ _03347_
+ sg13g2_a22oi_1
X_22936_ _03346_ _03347_ VPWR VGND _03348_ sg13g2_nand2_1
X_22937_ _08403_ _03348_ VPWR VGND _03349_ sg13g2_nand2_1
X_22938_ _03191_ _03321_ _03349_ VPWR VGND _03350_ sg13g2_nand3b_1
X_22939_ _03341_ _03345_ VPWR VGND _03351_ sg13g2_nand2_1
X_22940_ _00049_ VPWR VGND _03352_ sg13g2_inv_1
X_22941_ _03336_ _03338_ VPWR VGND _03353_ sg13g2_or2_1
X_22942_ _03353_ VPWR VGND _03354_ sg13g2_buf_2
X_22943_ _11132_ _00045_ VPWR VGND _03355_ sg13g2_nand2_1
X_22944_ _03293_ _03337_ _03355_ VPWR VGND _03356_ sg13g2_a21o_1
X_22945_ _03324_ _03329_ _03332_ VPWR VGND _03357_ sg13g2_a21o_1
X_22946_ _00047_ VPWR VGND _03358_ sg13g2_inv_1
X_22947_ _03334_ _03299_ _03358_ VPWR VGND _03359_ sg13g2_o21ai_1
X_22948_ _03249_ _03357_ _03359_ VPWR VGND _03360_ sg13g2_a21oi_1
X_22949_ _03356_ _03360_ _03277_ VPWR VGND _03361_ sg13g2_a21oi_1
X_22950_ _03301_ _03302_ VPWR VGND _03362_ sg13g2_or2_1
X_22951_ _03277_ _10957_ VPWR VGND _03363_ sg13g2_nand2_1
X_22952_ _03356_ _03360_ _03363_ VPWR VGND _03364_ sg13g2_a21oi_1
X_22953_ _03232_ _03354_ _03361_ _03362_ _03364_ VPWR 
+ VGND
+ _03365_ sg13g2_a221oi_1
X_22954_ _03365_ VPWR VGND _03366_ sg13g2_buf_2
X_22955_ _10794_ _03279_ _03280_ _03303_ VPWR VGND 
+ _03367_
+ sg13g2_nand4_1
X_22956_ _10795_ _10624_ VPWR VGND _03368_ sg13g2_nand2_1
X_22957_ _03352_ _03366_ _03367_ _03368_ VPWR VGND 
+ _03369_
+ sg13g2_a22oi_1
X_22958_ _03313_ _03351_ _03369_ VPWR VGND _03370_ sg13g2_a21oi_1
X_22959_ _03311_ _03313_ _03255_ _10794_ VPWR VGND 
+ _03371_
+ sg13g2_a22oi_1
X_22960_ _03003_ _03011_ VPWR VGND _03372_ sg13g2_nand2_1
X_22961_ _02969_ _02973_ VPWR VGND _03373_ sg13g2_nor2_1
X_22962_ _10458_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _03373_ _03202_ VPWR VGND 
+ _03374_
+ sg13g2_nor4_1
X_22963_ _03372_ _03208_ _03374_ VPWR VGND _03375_ sg13g2_nand3_1
X_22964_ _03016_ _03248_ _03322_ _03375_ VPWR VGND 
+ _03376_
+ sg13g2_or4_1
X_22965_ _03100_ _03112_ _03096_ _03053_ VPWR VGND 
+ _03377_
+ sg13g2_a22oi_1
X_22966_ _03305_ _03376_ _03377_ VPWR VGND _03378_ sg13g2_nor3_1
X_22967_ _09710_ _03371_ _03378_ VPWR VGND _03379_ sg13g2_o21ai_1
X_22968_ _03149_ _03348_ _03379_ VPWR VGND _03380_ sg13g2_or3_1
X_22969_ _03165_ _03170_ _03370_ _08403_ _03380_ VPWR 
+ VGND
+ _03381_ sg13g2_a221oi_1
X_22970_ _10624_ _03311_ VPWR VGND _03382_ sg13g2_nand2_1
X_22971_ _08980_ _03199_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ VPWR VGND _03383_ sg13g2_a21oi_1
X_22972_ _03104_ _03221_ _03225_ _03383_ VPWR VGND 
+ _03384_
+ sg13g2_nand4_1
X_22973_ _03156_ _03231_ _03253_ _03384_ VPWR VGND 
+ _03385_
+ sg13g2_nor4_1
X_22974_ _03159_ _03178_ _03382_ _03385_ VPWR VGND 
+ _03386_
+ sg13g2_nand4_1
X_22975_ _03311_ _03313_ VPWR VGND _03387_ sg13g2_nand2_1
X_22976_ _08403_ VPWR VGND _03388_ sg13g2_inv_1
X_22977_ _03387_ _03306_ _03388_ VPWR VGND _03389_ sg13g2_a21oi_1
X_22978_ _03188_ _03386_ _03389_ VPWR VGND _03390_ sg13g2_nor3_1
X_22979_ _03350_ _03381_ _03390_ VPWR VGND _03391_ sg13g2_o21ai_1
X_22980_ _03085_ _03168_ VPWR VGND _03392_ sg13g2_nand2_1
X_22981_ _09534_ _03084_ _03392_ VPWR VGND _03393_ sg13g2_a21oi_1
X_22982_ _03293_ _03337_ _03355_ VPWR VGND _03394_ sg13g2_a21oi_1
X_22983_ _03228_ _03333_ VPWR VGND _03395_ sg13g2_nor2_1
X_22984_ _03334_ _03299_ VPWR VGND _03396_ sg13g2_nor2_1
X_22985_ _10957_ _03394_ _03395_ _03396_ VPWR VGND 
+ _03397_
+ sg13g2_or4_1
X_22986_ _10957_ _03358_ _10960_ VPWR VGND _03398_ sg13g2_a21oi_1
X_22987_ _03277_ _03358_ VPWR VGND _03399_ sg13g2_nor2_1
X_22988_ _03397_ _03398_ _03399_ _03354_ VPWR VGND 
+ _03400_
+ sg13g2_a22oi_1
X_22989_ _10625_ _03400_ VPWR VGND _03401_ sg13g2_nand2_1
X_22990_ _10624_ _03352_ _10794_ VPWR VGND _03402_ sg13g2_a21oi_1
X_22991_ _03352_ _03366_ VPWR VGND _03403_ sg13g2_nor2_1
X_22992_ _03401_ _03402_ _03403_ _10794_ VPWR VGND 
+ _03404_
+ sg13g2_a22oi_1
X_22993_ _09914_ _09712_ _03017_ VPWR VGND _03405_ sg13g2_o21ai_1
X_22994_ _09914_ _03037_ _03405_ VPWR VGND _03406_ sg13g2_a21oi_1
X_22995_ _03285_ _03287_ _03289_ VPWR VGND _03407_ sg13g2_or3_1
X_22996_ _08980_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ VPWR VGND _03408_ sg13g2_nor2_1
X_22997_ _09150_ _03408_ _00040_ VPWR VGND _03409_ sg13g2_a21oi_1
X_22998_ _03024_ _03409_ VPWR VGND _03410_ sg13g2_nand2_1
X_22999_ _03062_ _03407_ _03396_ _03410_ VPWR VGND 
+ _03411_
+ sg13g2_or4_1
X_23000_ _03357_ _03394_ _03406_ _03411_ VPWR VGND 
+ _03412_
+ sg13g2_nor4_1
X_23001_ _03358_ _03232_ VPWR VGND _03413_ sg13g2_nor2_1
X_23002_ _03277_ _03354_ _03413_ VPWR VGND _03414_ sg13g2_o21ai_1
X_23003_ _03091_ _03404_ _03412_ _03414_ VPWR VGND 
+ _03415_
+ sg13g2_nand4_1
X_23004_ _03366_ _03313_ VPWR VGND _03416_ sg13g2_nor2b_1
X_23005_ _03341_ _03345_ _03400_ _03352_ _10795_ VPWR 
+ VGND
+ _03417_ sg13g2_a221oi_1
X_23006_ _03352_ _03400_ _03368_ VPWR VGND _03418_ sg13g2_a21oi_1
X_23007_ _03416_ _03417_ _03418_ VPWR VGND _03419_ sg13g2_nor3_1
X_23008_ _09709_ _08403_ _00050_ VPWR VGND _03420_ sg13g2_o21ai_1
X_23009_ _09709_ _03419_ _03420_ VPWR VGND _03421_ sg13g2_a21oi_1
X_23010_ _03393_ _03415_ _03421_ VPWR VGND _03422_ sg13g2_or3_1
X_23011_ _03422_ VPWR VGND _03423_ sg13g2_buf_1
X_23012_ _03341_ _03345_ VPWR VGND _03424_ sg13g2_and2_1
X_23013_ _03004_ _02980_ VPWR VGND _03425_ sg13g2_and2_1
X_23014_ _10455_ _02970_ _10621_ VPWR VGND _03426_ sg13g2_a21oi_1
X_23015_ _10458_ _03426_ _03194_ VPWR VGND _03427_ sg13g2_o21ai_1
X_23016_ _00044_ _03296_ _03425_ _03427_ VPWR VGND 
+ _03428_
+ sg13g2_nor4_1
X_23017_ _03047_ _03052_ _03275_ _03428_ VPWR VGND 
+ _03429_
+ sg13g2_nand4_1
X_23018_ _03057_ _03362_ _03429_ VPWR VGND _03430_ sg13g2_nor3_1
X_23019_ _03118_ _03424_ _03370_ _03430_ VPWR VGND 
+ _03431_
+ sg13g2_nand4_1
X_23020_ _00050_ VPWR VGND _03432_ sg13g2_inv_1
X_23021_ _09709_ _03346_ _03347_ VPWR VGND _03433_ sg13g2_nand3_1
X_23022_ _09710_ _08403_ VPWR VGND _03434_ sg13g2_nand2_1
X_23023_ _03432_ _03419_ _03433_ _03434_ VPWR VGND 
+ _03435_
+ sg13g2_a22oi_1
X_23024_ _03150_ _03431_ _03435_ VPWR VGND _03436_ sg13g2_nor3_1
X_23025_ _02978_ _02986_ _03198_ _03238_ _00042_ VPWR 
+ VGND
+ _03437_ sg13g2_a221oi_1
X_23026_ _02995_ _02965_ VPWR VGND _03438_ sg13g2_nor2_1
X_23027_ _10453_ _03044_ _03438_ VPWR VGND _03439_ sg13g2_o21ai_1
X_23028_ _03283_ _03437_ _03439_ VPWR VGND _03440_ sg13g2_nand3_1
X_23029_ _03037_ _03293_ _03337_ VPWR VGND _03441_ sg13g2_nand3_1
X_23030_ _03354_ _03440_ _03441_ VPWR VGND _03442_ sg13g2_nor3_1
X_23031_ _03080_ _03084_ _03366_ _03442_ VPWR VGND 
+ _03443_
+ sg13g2_nand4_1
X_23032_ _03086_ _03091_ _03118_ _09533_ _03092_ VPWR 
+ VGND
+ _03444_ sg13g2_a221oi_1
X_23033_ _03444_ _03419_ VPWR VGND _03445_ sg13g2_nand2b_1
X_23034_ _09709_ _08403_ VPWR VGND _03446_ sg13g2_nor2_1
X_23035_ _09709_ _03370_ _03404_ _03432_ _03446_ VPWR 
+ VGND
+ _03447_ sg13g2_a221oi_1
X_23036_ _03443_ _03445_ _03447_ VPWR VGND _03448_ sg13g2_nor3_1
X_23037_ _03436_ _03448_ VPWR VGND _03449_ sg13g2_nor2b_1
X_23038_ _03423_ _03449_ VPWR VGND _03450_ sg13g2_nor2_1
X_23039_ _03391_ _03450_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[0]\ sg13g2_xnor2_1
X_23040_ _03423_ _03449_ _03391_ VPWR VGND _03451_ sg13g2_o21ai_1
X_23041_ _03423_ _03448_ VPWR VGND _03452_ sg13g2_nand2b_1
X_23042_ _03183_ _03390_ _03321_ _03349_ VPWR VGND 
+ _03453_
+ sg13g2_nand4_1
X_23043_ _03453_ VPWR VGND _03454_ sg13g2_buf_1
X_23044_ _03452_ _03454_ VPWR VGND _03455_ sg13g2_xor2_1
X_23045_ _03451_ _03455_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[1]\ sg13g2_xnor2_1
X_23046_ _03452_ _03454_ VPWR VGND _03456_ sg13g2_nand2_1
X_23047_ _03452_ _03454_ VPWR VGND _03457_ sg13g2_nor2_1
X_23048_ _03451_ _03456_ _03457_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[2]\ sg13g2_a21oi_1
X_23049_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3028_q\ _07928_ VPWR VGND \atbs_core_0.adaptive_ctrl_0.n1658_o\ sg13g2_nand2b_1
X_23050_ \atbs_core_0.dac_control_0.n1942_q[0]\ _11609_ VPWR VGND \atbs_core_0.dac_control_0.n1904_o[0]\ sg13g2_nor2_1
X_23051_ \atbs_core_0.dac_control_0.n1942_q[1]\ \atbs_core_0.dac_control_0.n1942_q[0]\ VPWR VGND _03458_ sg13g2_xnor2_1
X_23052_ _11609_ _03458_ VPWR VGND \atbs_core_0.dac_control_0.n1904_o[1]\ sg13g2_nor2_1
X_23053_ _00058_ _11607_ VPWR VGND _03459_ sg13g2_xnor2_1
X_23054_ _11609_ _03459_ VPWR VGND \atbs_core_0.dac_control_0.n1904_o[2]\ sg13g2_nor2_1
X_23055_ \atbs_core_0.dac_control_1.n2091_q[0]\ _11834_ VPWR VGND \atbs_core_0.dac_control_1.n2053_o[0]\ sg13g2_nor2_1
X_23056_ \atbs_core_0.dac_control_1.n2091_q[1]\ \atbs_core_0.dac_control_1.n2091_q[0]\ VPWR VGND _03460_ sg13g2_xnor2_1
X_23057_ _11834_ _03460_ VPWR VGND \atbs_core_0.dac_control_1.n2053_o[1]\ sg13g2_nor2_1
X_23058_ _00059_ _11831_ VPWR VGND _03461_ sg13g2_xnor2_1
X_23059_ _11834_ _03461_ VPWR VGND \atbs_core_0.dac_control_1.n2053_o[2]\ sg13g2_nor2_1
X_23060_ \atbs_core_0.debouncer_0.bouncing_sync\ _11870_ VPWR VGND _03462_ sg13g2_xnor2_1
X_23061_ _11852_ _11851_ _03462_ VPWR VGND _03463_ sg13g2_nor3_1
X_23062_ _03463_ VPWR VGND _03464_ sg13g2_inv_1
X_23063_ _11869_ _03464_ VPWR VGND _03465_ sg13g2_nand2_1
X_23064_ _03465_ VPWR VGND _03466_ sg13g2_buf_1
X_23065_ _11855_ _03466_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[0]\ sg13g2_nor2_1
X_23066_ _11853_ _11862_ VPWR VGND _03467_ sg13g2_xnor2_1
X_23067_ _03466_ _03467_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[10]\ sg13g2_nor2_1
X_23068_ \atbs_core_0.debouncer_0.counter_value[11]\ _11863_ VPWR VGND _03468_ sg13g2_xnor2_1
X_23069_ _03466_ _03468_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[11]\ sg13g2_nor2_1
X_23070_ \atbs_core_0.debouncer_0.counter_value[12]\ _11865_ VPWR VGND _03469_ sg13g2_xnor2_1
X_23071_ _03463_ _03469_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[12]\ sg13g2_nor2_1
X_23072_ \atbs_core_0.debouncer_0.counter_value[12]\ _11865_ VPWR VGND _03470_ sg13g2_nand2_1
X_23073_ \atbs_core_0.debouncer_0.counter_value[13]\ _03470_ VPWR VGND _03471_ sg13g2_xor2_1
X_23074_ _03463_ _03471_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[13]\ sg13g2_nor2_1
X_23075_ \atbs_core_0.debouncer_0.counter_value[14]\ _11867_ VPWR VGND _03472_ sg13g2_xnor2_1
X_23076_ _03463_ _03472_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[14]\ sg13g2_nor2_1
X_23077_ \atbs_core_0.debouncer_0.counter_value[14]\ _11867_ VPWR VGND _03473_ sg13g2_nand2_1
X_23078_ \atbs_core_0.debouncer_0.counter_value[15]\ _03473_ VPWR VGND _03474_ sg13g2_xor2_1
X_23079_ _03463_ _03474_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[15]\ sg13g2_nor2_1
X_23080_ \atbs_core_0.debouncer_0.counter_value[1]\ _11855_ VPWR VGND _03475_ sg13g2_xnor2_1
X_23081_ _03466_ _03475_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[1]\ sg13g2_nor2_1
X_23082_ \atbs_core_0.debouncer_0.counter_value[1]\ _11855_ VPWR VGND _03476_ sg13g2_nand2_1
X_23083_ \atbs_core_0.debouncer_0.counter_value[2]\ _03476_ VPWR VGND _03477_ sg13g2_xor2_1
X_23084_ _03466_ _03477_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[2]\ sg13g2_nor2_1
X_23085_ _11854_ _11856_ VPWR VGND _03478_ sg13g2_xnor2_1
X_23086_ _03466_ _03478_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[3]\ sg13g2_nor2_1
X_23087_ \atbs_core_0.debouncer_0.counter_value[4]\ _11857_ VPWR VGND _03479_ sg13g2_xnor2_1
X_23088_ _03466_ _03479_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[4]\ sg13g2_nor2_1
X_23089_ \atbs_core_0.debouncer_0.counter_value[4]\ _11857_ VPWR VGND _03480_ sg13g2_nand2_1
X_23090_ \atbs_core_0.debouncer_0.counter_value[5]\ _03480_ VPWR VGND _03481_ sg13g2_xor2_1
X_23091_ _03466_ _03481_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[5]\ sg13g2_nor2_1
X_23092_ \atbs_core_0.debouncer_0.counter_value[6]\ _11859_ VPWR VGND _03482_ sg13g2_xnor2_1
X_23093_ _03466_ _03482_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[6]\ sg13g2_nor2_1
X_23094_ \atbs_core_0.debouncer_0.counter_value[6]\ _11859_ VPWR VGND _03483_ sg13g2_nand2_1
X_23095_ \atbs_core_0.debouncer_0.counter_value[7]\ _03483_ VPWR VGND _03484_ sg13g2_xor2_1
X_23096_ _03466_ _03484_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[7]\ sg13g2_nor2_1
X_23097_ \atbs_core_0.debouncer_0.counter_value[8]\ _11861_ VPWR VGND _03485_ sg13g2_xnor2_1
X_23098_ _03465_ _03485_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[8]\ sg13g2_nor2_1
X_23099_ \atbs_core_0.debouncer_0.counter_value[8]\ _11861_ VPWR VGND _03486_ sg13g2_nand2_1
X_23100_ \atbs_core_0.debouncer_0.counter_value[9]\ _03486_ VPWR VGND _03487_ sg13g2_xor2_1
X_23101_ _03465_ _03487_ VPWR VGND \atbs_core_0.debouncer_0.n1466_o[9]\ sg13g2_nor2_1
X_23102_ \atbs_core_0.debouncer_1.bouncing_sync\ _11898_ VPWR VGND _03488_ sg13g2_xnor2_1
X_23103_ _11880_ _11879_ _03488_ VPWR VGND _03489_ sg13g2_nor3_1
X_23104_ _03489_ VPWR VGND _03490_ sg13g2_inv_1
X_23105_ _11897_ _03490_ VPWR VGND _03491_ sg13g2_nand2_1
X_23106_ _03491_ VPWR VGND _03492_ sg13g2_buf_1
X_23107_ _11883_ _03492_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[0]\ sg13g2_nor2_1
X_23108_ _11881_ _11890_ VPWR VGND _03493_ sg13g2_xnor2_1
X_23109_ _03492_ _03493_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[10]\ sg13g2_nor2_1
X_23110_ \atbs_core_0.debouncer_1.counter_value[11]\ _11891_ VPWR VGND _03494_ sg13g2_xnor2_1
X_23111_ _03492_ _03494_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[11]\ sg13g2_nor2_1
X_23112_ \atbs_core_0.debouncer_1.counter_value[12]\ _11893_ VPWR VGND _03495_ sg13g2_xnor2_1
X_23113_ _03489_ _03495_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[12]\ sg13g2_nor2_1
X_23114_ \atbs_core_0.debouncer_1.counter_value[12]\ _11893_ VPWR VGND _03496_ sg13g2_nand2_1
X_23115_ \atbs_core_0.debouncer_1.counter_value[13]\ _03496_ VPWR VGND _03497_ sg13g2_xor2_1
X_23116_ _03489_ _03497_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[13]\ sg13g2_nor2_1
X_23117_ \atbs_core_0.debouncer_1.counter_value[14]\ _11895_ VPWR VGND _03498_ sg13g2_xnor2_1
X_23118_ _03489_ _03498_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[14]\ sg13g2_nor2_1
X_23119_ \atbs_core_0.debouncer_1.counter_value[14]\ _11895_ VPWR VGND _03499_ sg13g2_nand2_1
X_23120_ \atbs_core_0.debouncer_1.counter_value[15]\ _03499_ VPWR VGND _03500_ sg13g2_xor2_1
X_23121_ _03489_ _03500_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[15]\ sg13g2_nor2_1
X_23122_ \atbs_core_0.debouncer_1.counter_value[1]\ _11883_ VPWR VGND _03501_ sg13g2_xnor2_1
X_23123_ _03492_ _03501_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[1]\ sg13g2_nor2_1
X_23124_ \atbs_core_0.debouncer_1.counter_value[1]\ _11883_ VPWR VGND _03502_ sg13g2_nand2_1
X_23125_ \atbs_core_0.debouncer_1.counter_value[2]\ _03502_ VPWR VGND _03503_ sg13g2_xor2_1
X_23126_ _03492_ _03503_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[2]\ sg13g2_nor2_1
X_23127_ _11882_ _11884_ VPWR VGND _03504_ sg13g2_xnor2_1
X_23128_ _03492_ _03504_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[3]\ sg13g2_nor2_1
X_23129_ \atbs_core_0.debouncer_1.counter_value[4]\ _11885_ VPWR VGND _03505_ sg13g2_xnor2_1
X_23130_ _03492_ _03505_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[4]\ sg13g2_nor2_1
X_23131_ \atbs_core_0.debouncer_1.counter_value[4]\ _11885_ VPWR VGND _03506_ sg13g2_nand2_1
X_23132_ \atbs_core_0.debouncer_1.counter_value[5]\ _03506_ VPWR VGND _03507_ sg13g2_xor2_1
X_23133_ _03492_ _03507_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[5]\ sg13g2_nor2_1
X_23134_ \atbs_core_0.debouncer_1.counter_value[6]\ _11887_ VPWR VGND _03508_ sg13g2_xnor2_1
X_23135_ _03492_ _03508_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[6]\ sg13g2_nor2_1
X_23136_ \atbs_core_0.debouncer_1.counter_value[6]\ _11887_ VPWR VGND _03509_ sg13g2_nand2_1
X_23137_ \atbs_core_0.debouncer_1.counter_value[7]\ _03509_ VPWR VGND _03510_ sg13g2_xor2_1
X_23138_ _03492_ _03510_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[7]\ sg13g2_nor2_1
X_23139_ \atbs_core_0.debouncer_1.counter_value[8]\ _11889_ VPWR VGND _03511_ sg13g2_xnor2_1
X_23140_ _03491_ _03511_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[8]\ sg13g2_nor2_1
X_23141_ \atbs_core_0.debouncer_1.counter_value[8]\ _11889_ VPWR VGND _03512_ sg13g2_nand2_1
X_23142_ \atbs_core_0.debouncer_1.counter_value[9]\ _03512_ VPWR VGND _03513_ sg13g2_xor2_1
X_23143_ _03491_ _03513_ VPWR VGND \atbs_core_0.debouncer_1.n1466_o[9]\ sg13g2_nor2_1
X_23144_ \atbs_core_0.debouncer_2.bouncing_sync\ _11926_ VPWR VGND _03514_ sg13g2_xnor2_1
X_23145_ _11908_ _11907_ _03514_ VPWR VGND _03515_ sg13g2_nor3_1
X_23146_ _03515_ VPWR VGND _03516_ sg13g2_inv_1
X_23147_ _11925_ _03516_ VPWR VGND _03517_ sg13g2_nand2_1
X_23148_ _03517_ VPWR VGND _03518_ sg13g2_buf_1
X_23149_ _11911_ _03518_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[0]\ sg13g2_nor2_1
X_23150_ _11909_ _11918_ VPWR VGND _03519_ sg13g2_xnor2_1
X_23151_ _03518_ _03519_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[10]\ sg13g2_nor2_1
X_23152_ \atbs_core_0.debouncer_2.counter_value[11]\ _11919_ VPWR VGND _03520_ sg13g2_xnor2_1
X_23153_ _03518_ _03520_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[11]\ sg13g2_nor2_1
X_23154_ \atbs_core_0.debouncer_2.counter_value[12]\ _11921_ VPWR VGND _03521_ sg13g2_xnor2_1
X_23155_ _03515_ _03521_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[12]\ sg13g2_nor2_1
X_23156_ \atbs_core_0.debouncer_2.counter_value[12]\ _11921_ VPWR VGND _03522_ sg13g2_nand2_1
X_23157_ \atbs_core_0.debouncer_2.counter_value[13]\ _03522_ VPWR VGND _03523_ sg13g2_xor2_1
X_23158_ _03515_ _03523_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[13]\ sg13g2_nor2_1
X_23159_ \atbs_core_0.debouncer_2.counter_value[14]\ _11923_ VPWR VGND _03524_ sg13g2_xnor2_1
X_23160_ _03515_ _03524_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[14]\ sg13g2_nor2_1
X_23161_ \atbs_core_0.debouncer_2.counter_value[14]\ _11923_ VPWR VGND _03525_ sg13g2_nand2_1
X_23162_ \atbs_core_0.debouncer_2.counter_value[15]\ _03525_ VPWR VGND _03526_ sg13g2_xor2_1
X_23163_ _03515_ _03526_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[15]\ sg13g2_nor2_1
X_23164_ \atbs_core_0.debouncer_2.counter_value[1]\ _11911_ VPWR VGND _03527_ sg13g2_xnor2_1
X_23165_ _03518_ _03527_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[1]\ sg13g2_nor2_1
X_23166_ \atbs_core_0.debouncer_2.counter_value[1]\ _11911_ VPWR VGND _03528_ sg13g2_nand2_1
X_23167_ \atbs_core_0.debouncer_2.counter_value[2]\ _03528_ VPWR VGND _03529_ sg13g2_xor2_1
X_23168_ _03518_ _03529_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[2]\ sg13g2_nor2_1
X_23169_ _11910_ _11912_ VPWR VGND _03530_ sg13g2_xnor2_1
X_23170_ _03518_ _03530_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[3]\ sg13g2_nor2_1
X_23171_ \atbs_core_0.debouncer_2.counter_value[4]\ _11913_ VPWR VGND _03531_ sg13g2_xnor2_1
X_23172_ _03518_ _03531_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[4]\ sg13g2_nor2_1
X_23173_ \atbs_core_0.debouncer_2.counter_value[4]\ _11913_ VPWR VGND _03532_ sg13g2_nand2_1
X_23174_ \atbs_core_0.debouncer_2.counter_value[5]\ _03532_ VPWR VGND _03533_ sg13g2_xor2_1
X_23175_ _03518_ _03533_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[5]\ sg13g2_nor2_1
X_23176_ \atbs_core_0.debouncer_2.counter_value[6]\ _11915_ VPWR VGND _03534_ sg13g2_xnor2_1
X_23177_ _03518_ _03534_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[6]\ sg13g2_nor2_1
X_23178_ \atbs_core_0.debouncer_2.counter_value[6]\ _11915_ VPWR VGND _03535_ sg13g2_nand2_1
X_23179_ \atbs_core_0.debouncer_2.counter_value[7]\ _03535_ VPWR VGND _03536_ sg13g2_xor2_1
X_23180_ _03518_ _03536_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[7]\ sg13g2_nor2_1
X_23181_ \atbs_core_0.debouncer_2.counter_value[8]\ _11917_ VPWR VGND _03537_ sg13g2_xnor2_1
X_23182_ _03517_ _03537_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[8]\ sg13g2_nor2_1
X_23183_ \atbs_core_0.debouncer_2.counter_value[8]\ _11917_ VPWR VGND _03538_ sg13g2_nand2_1
X_23184_ \atbs_core_0.debouncer_2.counter_value[9]\ _03538_ VPWR VGND _03539_ sg13g2_xor2_1
X_23185_ _03517_ _03539_ VPWR VGND \atbs_core_0.debouncer_2.n1466_o[9]\ sg13g2_nor2_1
X_23186_ \atbs_core_0.debouncer_3.bouncing_sync\ _11953_ VPWR VGND _03540_ sg13g2_xnor2_1
X_23187_ _11936_ _11935_ _03540_ VPWR VGND _03541_ sg13g2_nor3_1
X_23188_ \atbs_core_0.debouncer_3.counter_value[15]\ _11951_ _03541_ VPWR VGND _03542_ sg13g2_a21o_1
X_23189_ _03542_ VPWR VGND _03543_ sg13g2_buf_1
X_23190_ _03543_ VPWR VGND _03544_ sg13g2_buf_1
X_23191_ _11941_ _03544_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[0]\ sg13g2_nor2_1
X_23192_ \atbs_core_0.debouncer_3.counter_value[9]\ _11947_ VPWR VGND _03545_ sg13g2_nand2_1
X_23193_ \atbs_core_0.debouncer_3.counter_value[10]\ _03545_ VPWR VGND _03546_ sg13g2_xor2_1
X_23194_ _03544_ _03546_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[10]\ sg13g2_nor2_1
X_23195_ _11938_ _11948_ VPWR VGND _03547_ sg13g2_xnor2_1
X_23196_ _03544_ _03547_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[11]\ sg13g2_nor2_1
X_23197_ \atbs_core_0.debouncer_3.counter_value[12]\ _11949_ VPWR VGND _03548_ sg13g2_xnor2_1
X_23198_ _03541_ _03548_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[12]\ sg13g2_nor2_1
X_23199_ \atbs_core_0.debouncer_3.counter_value[12]\ _11949_ VPWR VGND _03549_ sg13g2_nand2_1
X_23200_ \atbs_core_0.debouncer_3.counter_value[13]\ _03549_ VPWR VGND _03550_ sg13g2_xor2_1
X_23201_ _03541_ _03550_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[13]\ sg13g2_nor2_1
X_23202_ _11937_ _11950_ VPWR VGND _03551_ sg13g2_xnor2_1
X_23203_ _03541_ _03551_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[14]\ sg13g2_nor2_1
X_23204_ \atbs_core_0.debouncer_3.counter_value[15]\ _11951_ VPWR VGND _03552_ sg13g2_xnor2_1
X_23205_ _03541_ _03552_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[15]\ sg13g2_nor2_1
X_23206_ \atbs_core_0.debouncer_3.counter_value[1]\ _11941_ VPWR VGND _03553_ sg13g2_xnor2_1
X_23207_ _03544_ _03553_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[1]\ sg13g2_nor2_1
X_23208_ \atbs_core_0.debouncer_3.counter_value[1]\ _11941_ VPWR VGND _03554_ sg13g2_nand2_1
X_23209_ \atbs_core_0.debouncer_3.counter_value[2]\ _03554_ VPWR VGND _03555_ sg13g2_xor2_1
X_23210_ _03544_ _03555_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[2]\ sg13g2_nor2_1
X_23211_ _11940_ _11942_ VPWR VGND _03556_ sg13g2_xnor2_1
X_23212_ _03544_ _03556_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[3]\ sg13g2_nor2_1
X_23213_ \atbs_core_0.debouncer_3.counter_value[4]\ _11943_ VPWR VGND _03557_ sg13g2_xnor2_1
X_23214_ _03544_ _03557_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[4]\ sg13g2_nor2_1
X_23215_ \atbs_core_0.debouncer_3.counter_value[4]\ _11943_ VPWR VGND _03558_ sg13g2_nand2_1
X_23216_ \atbs_core_0.debouncer_3.counter_value[5]\ _03558_ VPWR VGND _03559_ sg13g2_xor2_1
X_23217_ _03544_ _03559_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[5]\ sg13g2_nor2_1
X_23218_ \atbs_core_0.debouncer_3.counter_value[6]\ _11945_ VPWR VGND _03560_ sg13g2_xnor2_1
X_23219_ _03544_ _03560_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[6]\ sg13g2_nor2_1
X_23220_ \atbs_core_0.debouncer_3.counter_value[6]\ _11945_ VPWR VGND _03561_ sg13g2_nand2_1
X_23221_ \atbs_core_0.debouncer_3.counter_value[7]\ _03561_ VPWR VGND _03562_ sg13g2_xor2_1
X_23222_ _03544_ _03562_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[7]\ sg13g2_nor2_1
X_23223_ _11939_ _11946_ VPWR VGND _03563_ sg13g2_xnor2_1
X_23224_ _03543_ _03563_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[8]\ sg13g2_nor2_1
X_23225_ \atbs_core_0.debouncer_3.counter_value[9]\ _11947_ VPWR VGND _03564_ sg13g2_xnor2_1
X_23226_ _03543_ _03564_ VPWR VGND \atbs_core_0.debouncer_3.n1466_o[9]\ sg13g2_nor2_1
X_23227_ \atbs_core_0.debouncer_4.bouncing_sync\ _11980_ VPWR VGND _03565_ sg13g2_xnor2_1
X_23228_ _11963_ _11962_ _03565_ VPWR VGND _03566_ sg13g2_nor3_1
X_23229_ \atbs_core_0.debouncer_4.counter_value[15]\ _11978_ _03566_ VPWR VGND _03567_ sg13g2_a21o_1
X_23230_ _03567_ VPWR VGND _03568_ sg13g2_buf_1
X_23231_ _03568_ VPWR VGND _03569_ sg13g2_buf_1
X_23232_ _11968_ _03569_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[0]\ sg13g2_nor2_1
X_23233_ \atbs_core_0.debouncer_4.counter_value[9]\ _11974_ VPWR VGND _03570_ sg13g2_nand2_1
X_23234_ \atbs_core_0.debouncer_4.counter_value[10]\ _03570_ VPWR VGND _03571_ sg13g2_xor2_1
X_23235_ _03569_ _03571_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[10]\ sg13g2_nor2_1
X_23236_ _11965_ _11975_ VPWR VGND _03572_ sg13g2_xnor2_1
X_23237_ _03569_ _03572_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[11]\ sg13g2_nor2_1
X_23238_ \atbs_core_0.debouncer_4.counter_value[12]\ _11976_ VPWR VGND _03573_ sg13g2_xnor2_1
X_23239_ _03566_ _03573_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[12]\ sg13g2_nor2_1
X_23240_ \atbs_core_0.debouncer_4.counter_value[12]\ _11976_ VPWR VGND _03574_ sg13g2_nand2_1
X_23241_ \atbs_core_0.debouncer_4.counter_value[13]\ _03574_ VPWR VGND _03575_ sg13g2_xor2_1
X_23242_ _03566_ _03575_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[13]\ sg13g2_nor2_1
X_23243_ _11964_ _11977_ VPWR VGND _03576_ sg13g2_xnor2_1
X_23244_ _03566_ _03576_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[14]\ sg13g2_nor2_1
X_23245_ \atbs_core_0.debouncer_4.counter_value[15]\ _11978_ VPWR VGND _03577_ sg13g2_xnor2_1
X_23246_ _03566_ _03577_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[15]\ sg13g2_nor2_1
X_23247_ \atbs_core_0.debouncer_4.counter_value[1]\ _11968_ VPWR VGND _03578_ sg13g2_xnor2_1
X_23248_ _03569_ _03578_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[1]\ sg13g2_nor2_1
X_23249_ \atbs_core_0.debouncer_4.counter_value[1]\ _11968_ VPWR VGND _03579_ sg13g2_nand2_1
X_23250_ \atbs_core_0.debouncer_4.counter_value[2]\ _03579_ VPWR VGND _03580_ sg13g2_xor2_1
X_23251_ _03569_ _03580_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[2]\ sg13g2_nor2_1
X_23252_ _11967_ _11969_ VPWR VGND _03581_ sg13g2_xnor2_1
X_23253_ _03569_ _03581_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[3]\ sg13g2_nor2_1
X_23254_ \atbs_core_0.debouncer_4.counter_value[4]\ _11970_ VPWR VGND _03582_ sg13g2_xnor2_1
X_23255_ _03569_ _03582_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[4]\ sg13g2_nor2_1
X_23256_ \atbs_core_0.debouncer_4.counter_value[4]\ _11970_ VPWR VGND _03583_ sg13g2_nand2_1
X_23257_ \atbs_core_0.debouncer_4.counter_value[5]\ _03583_ VPWR VGND _03584_ sg13g2_xor2_1
X_23258_ _03569_ _03584_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[5]\ sg13g2_nor2_1
X_23259_ \atbs_core_0.debouncer_4.counter_value[6]\ _11972_ VPWR VGND _03585_ sg13g2_xnor2_1
X_23260_ _03569_ _03585_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[6]\ sg13g2_nor2_1
X_23261_ \atbs_core_0.debouncer_4.counter_value[6]\ _11972_ VPWR VGND _03586_ sg13g2_nand2_1
X_23262_ \atbs_core_0.debouncer_4.counter_value[7]\ _03586_ VPWR VGND _03587_ sg13g2_xor2_1
X_23263_ _03569_ _03587_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[7]\ sg13g2_nor2_1
X_23264_ _11966_ _11973_ VPWR VGND _03588_ sg13g2_xnor2_1
X_23265_ _03568_ _03588_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[8]\ sg13g2_nor2_1
X_23266_ \atbs_core_0.debouncer_4.counter_value[9]\ _11974_ VPWR VGND _03589_ sg13g2_xnor2_1
X_23267_ _03568_ _03589_ VPWR VGND \atbs_core_0.debouncer_4.n1466_o[9]\ sg13g2_nor2_1
X_23268_ \atbs_core_0.debouncer_5.bouncing_sync\ _12008_ VPWR VGND _03590_ sg13g2_xnor2_1
X_23269_ _11989_ _11990_ _03590_ VPWR VGND _03591_ sg13g2_nor3_1
X_23270_ _03591_ VPWR VGND _03592_ sg13g2_inv_1
X_23271_ _12007_ _03592_ VPWR VGND _03593_ sg13g2_nand2_1
X_23272_ _03593_ VPWR VGND _03594_ sg13g2_buf_1
X_23273_ _11993_ _03594_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[0]\ sg13g2_nor2_1
X_23274_ _11991_ _12000_ VPWR VGND _03595_ sg13g2_xnor2_1
X_23275_ _03594_ _03595_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[10]\ sg13g2_nor2_1
X_23276_ \atbs_core_0.debouncer_5.counter_value[11]\ _12001_ VPWR VGND _03596_ sg13g2_xnor2_1
X_23277_ _03594_ _03596_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[11]\ sg13g2_nor2_1
X_23278_ \atbs_core_0.debouncer_5.counter_value[12]\ _12003_ VPWR VGND _03597_ sg13g2_xnor2_1
X_23279_ _03591_ _03597_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[12]\ sg13g2_nor2_1
X_23280_ \atbs_core_0.debouncer_5.counter_value[12]\ _12003_ VPWR VGND _03598_ sg13g2_nand2_1
X_23281_ \atbs_core_0.debouncer_5.counter_value[13]\ _03598_ VPWR VGND _03599_ sg13g2_xor2_1
X_23282_ _03591_ _03599_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[13]\ sg13g2_nor2_1
X_23283_ \atbs_core_0.debouncer_5.counter_value[14]\ _12005_ VPWR VGND _03600_ sg13g2_xnor2_1
X_23284_ _03591_ _03600_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[14]\ sg13g2_nor2_1
X_23285_ \atbs_core_0.debouncer_5.counter_value[14]\ _12005_ VPWR VGND _03601_ sg13g2_nand2_1
X_23286_ \atbs_core_0.debouncer_5.counter_value[15]\ _03601_ VPWR VGND _03602_ sg13g2_xor2_1
X_23287_ _03591_ _03602_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[15]\ sg13g2_nor2_1
X_23288_ \atbs_core_0.debouncer_5.counter_value[1]\ _11993_ VPWR VGND _03603_ sg13g2_xnor2_1
X_23289_ _03594_ _03603_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[1]\ sg13g2_nor2_1
X_23290_ \atbs_core_0.debouncer_5.counter_value[1]\ _11993_ VPWR VGND _03604_ sg13g2_nand2_1
X_23291_ \atbs_core_0.debouncer_5.counter_value[2]\ _03604_ VPWR VGND _03605_ sg13g2_xor2_1
X_23292_ _03594_ _03605_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[2]\ sg13g2_nor2_1
X_23293_ _11992_ _11994_ VPWR VGND _03606_ sg13g2_xnor2_1
X_23294_ _03594_ _03606_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[3]\ sg13g2_nor2_1
X_23295_ \atbs_core_0.debouncer_5.counter_value[4]\ _11995_ VPWR VGND _03607_ sg13g2_xnor2_1
X_23296_ _03594_ _03607_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[4]\ sg13g2_nor2_1
X_23297_ \atbs_core_0.debouncer_5.counter_value[4]\ _11995_ VPWR VGND _03608_ sg13g2_nand2_1
X_23298_ \atbs_core_0.debouncer_5.counter_value[5]\ _03608_ VPWR VGND _03609_ sg13g2_xor2_1
X_23299_ _03594_ _03609_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[5]\ sg13g2_nor2_1
X_23300_ \atbs_core_0.debouncer_5.counter_value[6]\ _11997_ VPWR VGND _03610_ sg13g2_xnor2_1
X_23301_ _03594_ _03610_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[6]\ sg13g2_nor2_1
X_23302_ \atbs_core_0.debouncer_5.counter_value[6]\ _11997_ VPWR VGND _03611_ sg13g2_nand2_1
X_23303_ \atbs_core_0.debouncer_5.counter_value[7]\ _03611_ VPWR VGND _03612_ sg13g2_xor2_1
X_23304_ _03594_ _03612_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[7]\ sg13g2_nor2_1
X_23305_ \atbs_core_0.debouncer_5.counter_value[8]\ _11999_ VPWR VGND _03613_ sg13g2_xnor2_1
X_23306_ _03593_ _03613_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[8]\ sg13g2_nor2_1
X_23307_ \atbs_core_0.debouncer_5.counter_value[8]\ _11999_ VPWR VGND _03614_ sg13g2_nand2_1
X_23308_ \atbs_core_0.debouncer_5.counter_value[9]\ _03614_ VPWR VGND _03615_ sg13g2_xor2_1
X_23309_ _03593_ _03615_ VPWR VGND \atbs_core_0.debouncer_5.n1466_o[9]\ sg13g2_nor2_1
X_23310_ _11423_ VPWR VGND _03616_ sg13g2_inv_1
X_23311_ _11438_ _02941_ _11421_ VPWR VGND _03617_ sg13g2_a21o_1
X_23312_ _11437_ _02941_ VPWR VGND _03618_ sg13g2_nand2_1
X_23313_ _03616_ _03617_ _03618_ _11421_ VPWR VGND 
+ _03619_
+ sg13g2_a22oi_1
X_23314_ _11416_ _02941_ _11444_ VPWR VGND _03620_ sg13g2_a21oi_1
X_23315_ _11444_ _03619_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ VPWR VGND _03621_ sg13g2_a21oi_1
X_23316_ _02942_ _03621_ VPWR VGND _03622_ sg13g2_nor2_1
X_23317_ _03619_ _03620_ _03622_ VPWR VGND _03623_ sg13g2_a21oi_1
X_23318_ _11375_ _11394_ _03623_ VPWR VGND _03624_ sg13g2_nor3_1
X_23319_ _11386_ _11375_ VPWR VGND _03625_ sg13g2_and2_1
X_23320_ _11386_ _11375_ VPWR VGND _03626_ sg13g2_nor2_1
X_23321_ _03625_ _03626_ _11395_ VPWR VGND _03627_ sg13g2_o21ai_1
X_23322_ _11394_ _03623_ _03627_ VPWR VGND _03628_ sg13g2_a21oi_1
X_23323_ _11386_ _03628_ _02941_ VPWR VGND _03629_ sg13g2_o21ai_1
X_23324_ _03624_ _03629_ VPWR VGND _03630_ sg13g2_nand2b_1
X_23325_ _11394_ _03623_ VPWR VGND _03631_ sg13g2_nor2_1
X_23326_ _03631_ _03625_ _03628_ VPWR VGND _03632_ sg13g2_a21oi_1
X_23327_ _11386_ _02941_ VPWR VGND _03633_ sg13g2_nand2_1
X_23328_ _11405_ _03633_ VPWR VGND _03634_ sg13g2_nor2_1
X_23329_ _11416_ _11486_ _02941_ VPWR VGND _03635_ sg13g2_nand3b_1
X_23330_ _11486_ _02941_ _03635_ VPWR VGND _03636_ sg13g2_o21ai_1
X_23331_ _11480_ _02942_ VPWR VGND _03637_ sg13g2_nor2_1
X_23332_ _03636_ _03637_ _11444_ VPWR VGND _03638_ sg13g2_mux2_1
X_23333_ _11421_ _11394_ VPWR VGND _03639_ sg13g2_nor2_1
X_23334_ _11423_ _11395_ _02941_ VPWR VGND _03640_ sg13g2_o21ai_1
X_23335_ _11395_ _11394_ VPWR VGND _03641_ sg13g2_xnor2_1
X_23336_ _11423_ _11421_ _03641_ VPWR VGND _03642_ sg13g2_nand3_1
X_23337_ _03616_ _11422_ _11395_ _11394_ VPWR VGND 
+ _03643_
+ sg13g2_nand4_1
X_23338_ _03642_ _03643_ VPWR VGND _03644_ sg13g2_nand2_1
X_23339_ _03639_ _03640_ _03644_ _02941_ VPWR VGND 
+ _03645_
+ sg13g2_a22oi_1
X_23340_ _11375_ _03633_ VPWR VGND _03646_ sg13g2_xnor2_1
X_23341_ _00085_ _00038_ _03645_ _03646_ VPWR VGND 
+ _03647_
+ sg13g2_nor4_1
X_23342_ _11410_ _11454_ VPWR VGND _03648_ sg13g2_nand2_1
X_23343_ _03632_ _03634_ _03638_ _03647_ _03648_ VPWR 
+ VGND
+ _03649_ sg13g2_a221oi_1
X_23344_ _11560_ _11455_ _00038_ _11533_ VPWR VGND 
+ _03650_
+ sg13g2_nor4_1
X_23345_ _11438_ _11552_ _11544_ VPWR VGND _03651_ sg13g2_nor3_1
X_23346_ _03630_ _03649_ _03650_ _03651_ VPWR VGND 
+ \atbs_core_0.n179_o\
+ sg13g2_a22oi_1
X_23347_ _11722_ _11629_ _11666_ _11683_ VPWR VGND 
+ _03652_
+ sg13g2_nor4_1
X_23348_ _11734_ _11730_ _11719_ VPWR VGND _03653_ sg13g2_nor3_1
X_23349_ _03652_ _03653_ VPWR VGND \atbs_core_0.n187_o\ sg13g2_nand2_1
X_23350_ _07657_ _07902_ VPWR VGND _03654_ sg13g2_nand2_1
X_23351_ _03654_ VPWR VGND _03655_ sg13g2_inv_1
X_23352_ _07909_ _03655_ _07917_ VPWR VGND _03656_ sg13g2_o21ai_1
X_23353_ _07709_ _12075_ VPWR VGND _03657_ sg13g2_nor2_1
X_23354_ \atbs_core_0.main_counter_value[7]\ VPWR VGND _03658_ sg13g2_inv_1
X_23355_ \atbs_core_0.main_counter_value[3]\ VPWR VGND _03659_ sg13g2_inv_1
X_23356_ _07700_ _07701_ \atbs_core_0.main_counter_value[2]\ VPWR VGND _03660_ sg13g2_nand3_1
X_23357_ _03659_ _03660_ VPWR VGND _03661_ sg13g2_nor2_1
X_23358_ _07697_ _07698_ \atbs_core_0.main_counter_value[6]\ _03661_ VPWR VGND 
+ _03662_
+ sg13g2_nand4_1
X_23359_ _03658_ _03662_ VPWR VGND _03663_ sg13g2_nor2_1
X_23360_ _07695_ \atbs_core_0.main_counter_value[19]\ VPWR VGND _03664_ sg13g2_nand2_1
X_23361_ \atbs_core_0.main_counter_value[13]\ _07692_ VPWR VGND _03665_ sg13g2_nand2_1
X_23362_ _07704_ _07705_ _03664_ _03665_ VPWR VGND 
+ _03666_
+ sg13g2_nor4_1
X_23363_ \atbs_core_0.main_counter_value[10]\ _07691_ _03663_ _03666_ VPWR VGND 
+ _03667_
+ sg13g2_nand4_1
X_23364_ _03656_ _03657_ _03667_ VPWR VGND _03668_ sg13g2_nand3_1
X_23365_ _03668_ VPWR VGND _03669_ sg13g2_buf_1
X_23366_ _03669_ VPWR VGND _03670_ sg13g2_buf_1
X_23367_ _07700_ _03670_ VPWR VGND \atbs_core_0.n268_o[0]\ sg13g2_nor2_1
X_23368_ \atbs_core_0.main_counter_value[10]\ VPWR VGND _03671_ sg13g2_inv_1
X_23369_ \atbs_core_0.main_counter_value[9]\ _07687_ _03663_ VPWR VGND _03672_ sg13g2_nand3_1
X_23370_ _03671_ _03672_ VPWR VGND _03673_ sg13g2_xnor2_1
X_23371_ _03670_ _03673_ VPWR VGND \atbs_core_0.n268_o[10]\ sg13g2_nor2_1
X_23372_ _03671_ _03672_ VPWR VGND _03674_ sg13g2_nor2_1
X_23373_ _07688_ _03674_ VPWR VGND _03675_ sg13g2_xnor2_1
X_23374_ _03670_ _03675_ VPWR VGND \atbs_core_0.n268_o[11]\ sg13g2_nor2_1
X_23375_ _07688_ _03674_ VPWR VGND _03676_ sg13g2_nand2_1
X_23376_ _07692_ _03676_ VPWR VGND _03677_ sg13g2_xor2_1
X_23377_ _03670_ _03677_ VPWR VGND \atbs_core_0.n268_o[12]\ sg13g2_nor2_1
X_23378_ _07688_ _07692_ _03674_ VPWR VGND _03678_ sg13g2_nand3_1
X_23379_ \atbs_core_0.main_counter_value[13]\ _03678_ VPWR VGND _03679_ sg13g2_xor2_1
X_23380_ _03670_ _03679_ VPWR VGND \atbs_core_0.n268_o[13]\ sg13g2_nor2_1
X_23381_ _03665_ _03676_ VPWR VGND _03680_ sg13g2_nor2_1
X_23382_ \atbs_core_0.main_counter_value[14]\ _03680_ VPWR VGND _03681_ sg13g2_xnor2_1
X_23383_ _03670_ _03681_ VPWR VGND \atbs_core_0.n268_o[14]\ sg13g2_nor2_1
X_23384_ \atbs_core_0.main_counter_value[14]\ _03680_ VPWR VGND _03682_ sg13g2_and2_1
X_23385_ _03682_ VPWR VGND _03683_ sg13g2_buf_1
X_23386_ _07689_ _03683_ VPWR VGND _03684_ sg13g2_xnor2_1
X_23387_ _03670_ _03684_ VPWR VGND \atbs_core_0.n268_o[15]\ sg13g2_nor2_1
X_23388_ _07689_ _03683_ VPWR VGND _03685_ sg13g2_nand2_1
X_23389_ _07705_ _03685_ VPWR VGND _03686_ sg13g2_xor2_1
X_23390_ _03670_ _03686_ VPWR VGND \atbs_core_0.n268_o[16]\ sg13g2_nor2_1
X_23391_ _07689_ _07705_ _03683_ VPWR VGND _03687_ sg13g2_and3_1
X_23392_ _03687_ VPWR VGND _03688_ sg13g2_buf_1
X_23393_ _07704_ _03688_ VPWR VGND _03689_ sg13g2_xnor2_1
X_23394_ _03670_ _03689_ VPWR VGND \atbs_core_0.n268_o[17]\ sg13g2_nor2_1
X_23395_ _07704_ _03688_ VPWR VGND _03690_ sg13g2_nand2_1
X_23396_ _07695_ _03690_ VPWR VGND _03691_ sg13g2_xor2_1
X_23397_ _03670_ _03691_ VPWR VGND \atbs_core_0.n268_o[18]\ sg13g2_nor2_1
X_23398_ _03669_ VPWR VGND _03692_ sg13g2_buf_1
X_23399_ _07704_ _07695_ _03688_ VPWR VGND _03693_ sg13g2_nand3_1
X_23400_ \atbs_core_0.main_counter_value[19]\ _03693_ VPWR VGND _03694_ sg13g2_xor2_1
X_23401_ _03692_ _03694_ VPWR VGND \atbs_core_0.n268_o[19]\ sg13g2_nor2_1
X_23402_ _07700_ _07701_ VPWR VGND _03695_ sg13g2_xnor2_1
X_23403_ _03692_ _03695_ VPWR VGND \atbs_core_0.n268_o[1]\ sg13g2_nor2_1
X_23404_ _07700_ _07701_ VPWR VGND _03696_ sg13g2_nand2_1
X_23405_ \atbs_core_0.main_counter_value[2]\ _03696_ VPWR VGND _03697_ sg13g2_xor2_1
X_23406_ _03692_ _03697_ VPWR VGND \atbs_core_0.n268_o[2]\ sg13g2_nor2_1
X_23407_ _03659_ _03660_ VPWR VGND _03698_ sg13g2_xnor2_1
X_23408_ _03692_ _03698_ VPWR VGND \atbs_core_0.n268_o[3]\ sg13g2_nor2_1
X_23409_ _07698_ _03661_ VPWR VGND _03699_ sg13g2_xnor2_1
X_23410_ _03692_ _03699_ VPWR VGND \atbs_core_0.n268_o[4]\ sg13g2_nor2_1
X_23411_ _07698_ _03661_ VPWR VGND _03700_ sg13g2_nand2_1
X_23412_ _07697_ _03700_ VPWR VGND _03701_ sg13g2_xor2_1
X_23413_ _03692_ _03701_ VPWR VGND \atbs_core_0.n268_o[5]\ sg13g2_nor2_1
X_23414_ _07697_ _07698_ _03661_ VPWR VGND _03702_ sg13g2_nand3_1
X_23415_ \atbs_core_0.main_counter_value[6]\ _03702_ VPWR VGND _03703_ sg13g2_xor2_1
X_23416_ _03692_ _03703_ VPWR VGND \atbs_core_0.n268_o[6]\ sg13g2_nor2_1
X_23417_ _03658_ _03662_ VPWR VGND _03704_ sg13g2_xnor2_1
X_23418_ _03692_ _03704_ VPWR VGND \atbs_core_0.n268_o[7]\ sg13g2_nor2_1
X_23419_ _07687_ _03663_ VPWR VGND _03705_ sg13g2_xnor2_1
X_23420_ _03692_ _03705_ VPWR VGND \atbs_core_0.n268_o[8]\ sg13g2_nor2_1
X_23421_ _07687_ _03663_ VPWR VGND _03706_ sg13g2_nand2_1
X_23422_ \atbs_core_0.main_counter_value[9]\ _03706_ VPWR VGND _03707_ sg13g2_xor2_1
X_23423_ _03692_ _03707_ VPWR VGND \atbs_core_0.n268_o[9]\ sg13g2_nor2_1
X_23424_ _07903_ _03654_ VPWR VGND _03708_ sg13g2_nand2_1
X_23425_ _07905_ _02951_ VPWR VGND _03709_ sg13g2_nor2b_1
X_23426_ _08009_ _03708_ _03709_ VPWR VGND _03710_ sg13g2_a21oi_1
X_23427_ _07903_ _02946_ VPWR VGND _03711_ sg13g2_nand2_1
X_23428_ _07909_ _03711_ VPWR VGND _03712_ sg13g2_nand2_1
X_23429_ _07905_ _03712_ _07684_ VPWR VGND _03713_ sg13g2_a21o_1
X_23430_ _07682_ _03710_ _03713_ VPWR VGND \atbs_core_0.n453_o[1]\ sg13g2_o21ai_1
X_23431_ _07684_ _03711_ _07915_ VPWR VGND _03714_ sg13g2_o21ai_1
X_23432_ _07905_ _03654_ VPWR VGND _03715_ sg13g2_nand2_1
X_23433_ _08009_ _03714_ _03715_ _07681_ VPWR VGND 
+ _03716_
+ sg13g2_a22oi_1
X_23434_ _03716_ VPWR VGND \atbs_core_0.n453_o[2]\ sg13g2_inv_1
X_23435_ _07921_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ VPWR VGND \atbs_core_0.spike_encoder_0.n2244_o\ sg13g2_and2_1
X_23436_ _07921_ _07733_ VPWR VGND \atbs_core_0.spike_encoder_0.n2250_o\ sg13g2_and2_1
X_23437_ _07541_ VPWR VGND _03717_ sg13g2_buf_1
X_23438_ _03717_ VPWR VGND _03718_ sg13g2_buf_1
X_23439_ _03718_ VPWR VGND _03719_ sg13g2_buf_1
X_23440_ _07547_ VPWR VGND _03720_ sg13g2_buf_1
X_23441_ _03720_ VPWR VGND _03721_ sg13g2_buf_1
X_23442_ _07552_ VPWR VGND _03722_ sg13g2_buf_1
X_23443_ _03722_ VPWR VGND _03723_ sg13g2_buf_1
X_23444_ _03723_ VPWR VGND _03724_ sg13g2_buf_1
X_23445_ _03724_ VPWR VGND _03725_ sg13g2_buf_1
X_23446_ _12091_ VPWR VGND _03726_ sg13g2_buf_1
X_23447_ _03726_ VPWR VGND _03727_ sg13g2_buf_1
X_23448_ _03727_ VPWR VGND _03728_ sg13g2_buf_1
X_23449_ _03728_ VPWR VGND _03729_ sg13g2_buf_1
X_23450_ _12080_ VPWR VGND _03730_ sg13g2_buf_1
X_23451_ _07528_ _03730_ _07560_ VPWR VGND _03731_ sg13g2_nor3_1
X_23452_ _03731_ VPWR VGND _03732_ sg13g2_buf_1
X_23453_ _03732_ VPWR VGND _03733_ sg13g2_buf_1
X_23454_ _12081_ _12082_ VPWR VGND _03734_ sg13g2_nand2_1
X_23455_ _03734_ VPWR VGND _03735_ sg13g2_buf_1
X_23456_ _03735_ VPWR VGND _03736_ sg13g2_buf_1
X_23457_ _03736_ VPWR VGND _03737_ sg13g2_buf_1
X_23458_ _02698_ VPWR VGND _03738_ sg13g2_buf_1
X_23459_ _03738_ VPWR VGND _03739_ sg13g2_buf_1
X_23460_ _03739_ VPWR VGND _03740_ sg13g2_buf_1
X_23461_ _07558_ VPWR VGND _03741_ sg13g2_buf_1
X_23462_ _03741_ VPWR VGND _03742_ sg13g2_buf_2
X_23463_ _03742_ VPWR VGND _03743_ sg13g2_buf_1
X_23464_ _03743_ VPWR VGND _03744_ sg13g2_buf_1
X_23465_ _02709_ VPWR VGND _03745_ sg13g2_buf_1
X_23466_ _03745_ VPWR VGND _03746_ sg13g2_buf_1
X_23467_ _03746_ VPWR VGND _03747_ sg13g2_buf_1
X_23468_ _03747_ _02391_ VPWR VGND _03748_ sg13g2_nor2_1
X_23469_ _07558_ VPWR VGND _03749_ sg13g2_buf_1
X_23470_ _03749_ VPWR VGND _03750_ sg13g2_buf_1
X_23471_ _03750_ VPWR VGND _03751_ sg13g2_buf_1
X_23472_ _02411_ _03751_ VPWR VGND _03752_ sg13g2_nor2_1
X_23473_ _02710_ VPWR VGND _03753_ sg13g2_buf_1
X_23474_ _03753_ VPWR VGND _03754_ sg13g2_buf_1
X_23475_ _03754_ VPWR VGND _03755_ sg13g2_buf_1
X_23476_ _03744_ _03748_ _03752_ _03755_ VPWR VGND 
+ _03756_
+ sg13g2_a22oi_1
X_23477_ _03730_ VPWR VGND _03757_ sg13g2_buf_1
X_23478_ _03757_ VPWR VGND _03758_ sg13g2_buf_1
X_23479_ _03758_ VPWR VGND _03759_ sg13g2_buf_1
X_23480_ _02710_ VPWR VGND _03760_ sg13g2_buf_1
X_23481_ _03760_ VPWR VGND _03761_ sg13g2_buf_1
X_23482_ _07526_ VPWR VGND _03762_ sg13g2_buf_1
X_23483_ _03762_ VPWR VGND _03763_ sg13g2_buf_1
X_23484_ _03763_ VPWR VGND _03764_ sg13g2_buf_1
X_23485_ _02391_ _03764_ VPWR VGND _03765_ sg13g2_nand2b_1
X_23486_ _03761_ _02411_ _03765_ VPWR VGND _03766_ sg13g2_o21ai_1
X_23487_ _02698_ VPWR VGND _03767_ sg13g2_buf_1
X_23488_ _03767_ VPWR VGND _03768_ sg13g2_buf_1
X_23489_ _03768_ VPWR VGND _03769_ sg13g2_buf_1
X_23490_ _03759_ _03766_ _03769_ VPWR VGND _03770_ sg13g2_a21oi_1
X_23491_ _03740_ _03756_ _03770_ VPWR VGND _03771_ sg13g2_a21oi_1
X_23492_ _00111_ _03733_ _03737_ _02430_ _03771_ VPWR 
+ VGND
+ _03772_ sg13g2_a221oi_1
X_23493_ _03726_ VPWR VGND _03773_ sg13g2_buf_1
X_23494_ _03773_ VPWR VGND _03774_ sg13g2_buf_1
X_23495_ _03774_ VPWR VGND _03775_ sg13g2_buf_1
X_23496_ _12085_ VPWR VGND _03776_ sg13g2_buf_1
X_23497_ \atbs_core_0.spike_memory_0.n2401_o[0]\ _03776_ VPWR VGND _03777_ sg13g2_nor2_1
X_23498_ _07563_ VPWR VGND _03778_ sg13g2_buf_1
X_23499_ _03778_ VPWR VGND _03779_ sg13g2_buf_1
X_23500_ _07552_ VPWR VGND _03780_ sg13g2_buf_1
X_23501_ \atbs_core_0.spike_memory_0.n2398_o[0]\ _03779_ _03780_ VPWR VGND _03781_ sg13g2_o21ai_1
X_23502_ _03742_ VPWR VGND _03782_ sg13g2_buf_1
X_23503_ _02711_ _02523_ VPWR VGND _03783_ sg13g2_nor2_1
X_23504_ _07558_ VPWR VGND _03784_ sg13g2_buf_1
X_23505_ _03784_ VPWR VGND _03785_ sg13g2_buf_1
X_23506_ _02544_ _03785_ VPWR VGND _03786_ sg13g2_nor2_1
X_23507_ _03745_ VPWR VGND _03787_ sg13g2_buf_1
X_23508_ _03787_ VPWR VGND _03788_ sg13g2_buf_1
X_23509_ _03782_ _03783_ _03786_ _03788_ VPWR VGND 
+ _03789_
+ sg13g2_a22oi_1
X_23510_ _03757_ VPWR VGND _03790_ sg13g2_buf_1
X_23511_ _03762_ VPWR VGND _03791_ sg13g2_buf_1
X_23512_ _02523_ _03791_ VPWR VGND _03792_ sg13g2_nand2b_1
X_23513_ _03746_ _02544_ _03792_ VPWR VGND _03793_ sg13g2_o21ai_1
X_23514_ _03790_ _03793_ _03768_ VPWR VGND _03794_ sg13g2_a21oi_1
X_23515_ _02700_ _03789_ _03794_ VPWR VGND _03795_ sg13g2_a21oi_1
X_23516_ _03777_ _03781_ _03795_ VPWR VGND _03796_ sg13g2_or3_1
X_23517_ _03775_ _03796_ VPWR VGND _03797_ sg13g2_nand2_1
X_23518_ _03729_ _03772_ _03797_ VPWR VGND _03798_ sg13g2_o21ai_1
X_23519_ _12090_ _07555_ VPWR VGND _03799_ sg13g2_nand2_1
X_23520_ _03799_ VPWR VGND _03800_ sg13g2_buf_1
X_23521_ _03800_ VPWR VGND _03801_ sg13g2_buf_1
X_23522_ _12084_ VPWR VGND _03802_ sg13g2_buf_1
X_23523_ _03802_ VPWR VGND _03803_ sg13g2_buf_1
X_23524_ _03803_ VPWR VGND _03804_ sg13g2_buf_1
X_23525_ \atbs_core_0.spike_memory_0.n2397_o[0]\ _03804_ VPWR VGND _03805_ sg13g2_nor2_1
X_23526_ _03778_ VPWR VGND _03806_ sg13g2_buf_1
X_23527_ _03806_ VPWR VGND _03807_ sg13g2_buf_1
X_23528_ \atbs_core_0.spike_memory_0.n2394_o[0]\ _03807_ VPWR VGND _03808_ sg13g2_nor2_1
X_23529_ _07525_ VPWR VGND _03809_ sg13g2_buf_1
X_23530_ _03809_ VPWR VGND _03810_ sg13g2_buf_1
X_23531_ _03810_ VPWR VGND _03811_ sg13g2_buf_1
X_23532_ _03811_ VPWR VGND _03812_ sg13g2_buf_1
X_23533_ _03742_ VPWR VGND _03813_ sg13g2_buf_1
X_23534_ _03813_ VPWR VGND _03814_ sg13g2_buf_1
X_23535_ _03745_ VPWR VGND _03815_ sg13g2_buf_1
X_23536_ _03815_ VPWR VGND _03816_ sg13g2_buf_1
X_23537_ _03816_ _02475_ VPWR VGND _03817_ sg13g2_nor2_1
X_23538_ _03784_ VPWR VGND _03818_ sg13g2_buf_1
X_23539_ _03818_ VPWR VGND _03819_ sg13g2_buf_1
X_23540_ _02497_ _03819_ VPWR VGND _03820_ sg13g2_nor2_1
X_23541_ _03745_ VPWR VGND _03821_ sg13g2_buf_1
X_23542_ _03821_ VPWR VGND _03822_ sg13g2_buf_1
X_23543_ _03822_ VPWR VGND _03823_ sg13g2_buf_1
X_23544_ _03814_ _03817_ _03820_ _03823_ VPWR VGND 
+ _03824_
+ sg13g2_a22oi_1
X_23545_ _03790_ VPWR VGND _03825_ sg13g2_buf_1
X_23546_ _03821_ VPWR VGND _03826_ sg13g2_buf_1
X_23547_ _03791_ VPWR VGND _03827_ sg13g2_buf_1
X_23548_ _02475_ _03827_ VPWR VGND _03828_ sg13g2_nand2b_1
X_23549_ _03826_ _02497_ _03828_ VPWR VGND _03829_ sg13g2_o21ai_1
X_23550_ _03767_ VPWR VGND _03830_ sg13g2_buf_1
X_23551_ _03830_ VPWR VGND _03831_ sg13g2_buf_1
X_23552_ _03825_ _03829_ _03831_ VPWR VGND _03832_ sg13g2_a21oi_1
X_23553_ _03812_ _03824_ _03832_ VPWR VGND _03833_ sg13g2_a21oi_1
X_23554_ _03805_ _03808_ _03833_ VPWR VGND _03834_ sg13g2_nor3_1
X_23555_ _03778_ VPWR VGND _03835_ sg13g2_buf_1
X_23556_ _03835_ VPWR VGND _03836_ sg13g2_buf_1
X_23557_ \atbs_core_0.spike_memory_0.n2405_o[0]\ _03736_ VPWR VGND _03837_ sg13g2_nand2b_1
X_23558_ \atbs_core_0.spike_memory_0.n2402_o[0]\ _03836_ _03837_ VPWR VGND _03838_ sg13g2_o21ai_1
X_23559_ _03767_ VPWR VGND _03839_ sg13g2_buf_1
X_23560_ _03839_ VPWR VGND _03840_ sg13g2_buf_1
X_23561_ _03840_ VPWR VGND _03841_ sg13g2_buf_1
X_23562_ _03749_ VPWR VGND _03842_ sg13g2_buf_1
X_23563_ _03842_ VPWR VGND _03843_ sg13g2_buf_1
X_23564_ _03843_ VPWR VGND _03844_ sg13g2_buf_1
X_23565_ _07526_ VPWR VGND _03845_ sg13g2_buf_1
X_23566_ _03845_ VPWR VGND _03846_ sg13g2_buf_1
X_23567_ _03846_ VPWR VGND _03847_ sg13g2_buf_1
X_23568_ _03847_ VPWR VGND _03848_ sg13g2_buf_1
X_23569_ _03848_ _02570_ VPWR VGND _03849_ sg13g2_nor2_1
X_23570_ _07558_ VPWR VGND _03850_ sg13g2_buf_1
X_23571_ _03850_ VPWR VGND _03851_ sg13g2_buf_1
X_23572_ _03851_ VPWR VGND _03852_ sg13g2_buf_1
X_23573_ _02592_ _03852_ VPWR VGND _03853_ sg13g2_nor2_1
X_23574_ _03845_ VPWR VGND _03854_ sg13g2_buf_1
X_23575_ _03854_ VPWR VGND _03855_ sg13g2_buf_1
X_23576_ _03855_ VPWR VGND _03856_ sg13g2_buf_1
X_23577_ _03856_ VPWR VGND _03857_ sg13g2_buf_1
X_23578_ _03844_ _03849_ _03853_ _03857_ VPWR VGND 
+ _03858_
+ sg13g2_a22oi_1
X_23579_ _03730_ VPWR VGND _03859_ sg13g2_buf_1
X_23580_ _03859_ VPWR VGND _03860_ sg13g2_buf_1
X_23581_ _03860_ VPWR VGND _03861_ sg13g2_buf_1
X_23582_ _02709_ VPWR VGND _03862_ sg13g2_buf_1
X_23583_ _03862_ VPWR VGND _03863_ sg13g2_buf_1
X_23584_ _03863_ VPWR VGND _03864_ sg13g2_buf_1
X_23585_ _02570_ _03864_ VPWR VGND _03865_ sg13g2_nand2b_1
X_23586_ _03856_ _02592_ _03865_ VPWR VGND _03866_ sg13g2_o21ai_1
X_23587_ _02698_ VPWR VGND _03867_ sg13g2_buf_1
X_23588_ _03867_ VPWR VGND _03868_ sg13g2_buf_1
X_23589_ _03868_ VPWR VGND _03869_ sg13g2_buf_1
X_23590_ _03861_ _03866_ _03869_ VPWR VGND _03870_ sg13g2_a21oi_1
X_23591_ _03841_ _03858_ _03870_ VPWR VGND _03871_ sg13g2_a21oi_1
X_23592_ _03774_ VPWR VGND _03872_ sg13g2_buf_1
X_23593_ _03838_ _03871_ _03872_ VPWR VGND _03873_ sg13g2_o21ai_1
X_23594_ _03801_ _03834_ _03873_ VPWR VGND _03874_ sg13g2_o21ai_1
X_23595_ _03725_ _03798_ _03874_ _03796_ VPWR VGND 
+ _03875_
+ sg13g2_a22oi_1
X_23596_ _12085_ VPWR VGND _03876_ sg13g2_buf_1
X_23597_ _03876_ VPWR VGND _03877_ sg13g2_buf_1
X_23598_ \atbs_core_0.spike_memory_0.n2365_o[0]\ _03877_ VPWR VGND _03878_ sg13g2_nor2_1
X_23599_ \atbs_core_0.spike_memory_0.n2362_o[0]\ _03836_ VPWR VGND _03879_ sg13g2_nor2_1
X_23600_ _02700_ VPWR VGND _03880_ sg13g2_buf_1
X_23601_ _03782_ VPWR VGND _03881_ sg13g2_buf_1
X_23602_ _02711_ VPWR VGND _03882_ sg13g2_buf_1
X_23603_ _03882_ _12625_ VPWR VGND _03883_ sg13g2_nor2_1
X_23604_ _03818_ VPWR VGND _03884_ sg13g2_buf_1
X_23605_ _12624_ _03884_ VPWR VGND _03885_ sg13g2_nor2_1
X_23606_ _02711_ VPWR VGND _03886_ sg13g2_buf_1
X_23607_ _03886_ VPWR VGND _03887_ sg13g2_buf_1
X_23608_ _03881_ _03883_ _03885_ _03887_ VPWR VGND 
+ _03888_
+ sg13g2_a22oi_1
X_23609_ _03790_ VPWR VGND _03889_ sg13g2_buf_1
X_23610_ _07526_ VPWR VGND _03890_ sg13g2_buf_1
X_23611_ _03890_ VPWR VGND _03891_ sg13g2_buf_1
X_23612_ _03891_ VPWR VGND _03892_ sg13g2_buf_1
X_23613_ _12625_ _03892_ VPWR VGND _03893_ sg13g2_nand2b_1
X_23614_ _03886_ _12624_ _03893_ VPWR VGND _03894_ sg13g2_o21ai_1
X_23615_ _03768_ VPWR VGND _03895_ sg13g2_buf_1
X_23616_ _03889_ _03894_ _03895_ VPWR VGND _03896_ sg13g2_a21oi_1
X_23617_ _03880_ _03888_ _03896_ VPWR VGND _03897_ sg13g2_a21oi_1
X_23618_ _03728_ _03878_ _03879_ _03897_ VPWR VGND 
+ _03898_
+ sg13g2_nor4_1
X_23619_ _07555_ VPWR VGND _03899_ sg13g2_buf_1
X_23620_ _03899_ VPWR VGND _03900_ sg13g2_buf_1
X_23621_ _03776_ VPWR VGND _03901_ sg13g2_buf_1
X_23622_ \atbs_core_0.spike_memory_0.n2373_o[0]\ _03901_ VPWR VGND _03902_ sg13g2_nor2_1
X_23623_ _03835_ VPWR VGND _03903_ sg13g2_buf_1
X_23624_ \atbs_core_0.spike_memory_0.n2370_o[0]\ _03903_ VPWR VGND _03904_ sg13g2_nor2_1
X_23625_ _03811_ VPWR VGND _03905_ sg13g2_buf_1
X_23626_ _03813_ VPWR VGND _03906_ sg13g2_buf_1
X_23627_ _03821_ VPWR VGND _03907_ sg13g2_buf_1
X_23628_ _03907_ _02079_ VPWR VGND _03908_ sg13g2_nor2_1
X_23629_ _03818_ VPWR VGND _03909_ sg13g2_buf_1
X_23630_ _02102_ _03909_ VPWR VGND _03910_ sg13g2_nor2_1
X_23631_ _03826_ VPWR VGND _03911_ sg13g2_buf_1
X_23632_ _03906_ _03908_ _03910_ _03911_ VPWR VGND 
+ _03912_
+ sg13g2_a22oi_1
X_23633_ _03790_ VPWR VGND _03913_ sg13g2_buf_1
X_23634_ _02711_ VPWR VGND _03914_ sg13g2_buf_1
X_23635_ _03890_ VPWR VGND _03915_ sg13g2_buf_1
X_23636_ _03915_ VPWR VGND _03916_ sg13g2_buf_1
X_23637_ _02079_ _03916_ VPWR VGND _03917_ sg13g2_nand2b_1
X_23638_ _03914_ _02102_ _03917_ VPWR VGND _03918_ sg13g2_o21ai_1
X_23639_ _03830_ VPWR VGND _03919_ sg13g2_buf_1
X_23640_ _03913_ _03918_ _03919_ VPWR VGND _03920_ sg13g2_a21oi_1
X_23641_ _03905_ _03912_ _03920_ VPWR VGND _03921_ sg13g2_a21oi_1
X_23642_ _03900_ _03902_ _03904_ _03921_ VPWR VGND 
+ _03922_
+ sg13g2_nor4_1
X_23643_ _03724_ _03898_ _03922_ VPWR VGND _03923_ sg13g2_nor3_1
X_23644_ _12090_ VPWR VGND _03924_ sg13g2_buf_1
X_23645_ _03924_ VPWR VGND _03925_ sg13g2_buf_1
X_23646_ _03727_ VPWR VGND _03926_ sg13g2_buf_1
X_23647_ \atbs_core_0.spike_memory_0.n2361_o[0]\ _12087_ VPWR VGND _03927_ sg13g2_nor2_1
X_23648_ \atbs_core_0.spike_memory_0.n2358_o[0]\ _03903_ VPWR VGND _03928_ sg13g2_nor2_1
X_23649_ _03813_ VPWR VGND _03929_ sg13g2_buf_1
X_23650_ _03821_ VPWR VGND _03930_ sg13g2_buf_1
X_23651_ _03930_ _02057_ VPWR VGND _03931_ sg13g2_nor2_1
X_23652_ _03818_ VPWR VGND _03932_ sg13g2_buf_1
X_23653_ _02229_ _03932_ VPWR VGND _03933_ sg13g2_nor2_1
X_23654_ _03914_ VPWR VGND _03934_ sg13g2_buf_1
X_23655_ _03929_ _03931_ _03933_ _03934_ VPWR VGND 
+ _03935_
+ sg13g2_a22oi_1
X_23656_ _03790_ VPWR VGND _03936_ sg13g2_buf_1
X_23657_ _03791_ VPWR VGND _03937_ sg13g2_buf_1
X_23658_ _02057_ _03937_ VPWR VGND _03938_ sg13g2_nand2b_1
X_23659_ _02712_ _02229_ _03938_ VPWR VGND _03939_ sg13g2_o21ai_1
X_23660_ _03768_ VPWR VGND _03940_ sg13g2_buf_1
X_23661_ _03936_ _03939_ _03940_ VPWR VGND _03941_ sg13g2_a21oi_1
X_23662_ _02701_ _03935_ _03941_ VPWR VGND _03942_ sg13g2_a21oi_1
X_23663_ _03926_ _03927_ _03928_ _03942_ VPWR VGND 
+ _03943_
+ sg13g2_nor4_1
X_23664_ _03776_ VPWR VGND _03944_ sg13g2_buf_1
X_23665_ \atbs_core_0.spike_memory_0.n2369_o[0]\ _03944_ VPWR VGND _03945_ sg13g2_nor2_1
X_23666_ _03806_ VPWR VGND _03946_ sg13g2_buf_1
X_23667_ \atbs_core_0.spike_memory_0.n2366_o[0]\ _03946_ VPWR VGND _03947_ sg13g2_nor2_1
X_23668_ _03811_ VPWR VGND _03948_ sg13g2_buf_1
X_23669_ _03855_ VPWR VGND _03949_ sg13g2_buf_1
X_23670_ _03949_ _02024_ VPWR VGND _03950_ sg13g2_nor2_1
X_23671_ _03784_ VPWR VGND _03951_ sg13g2_buf_1
X_23672_ _03951_ VPWR VGND _03952_ sg13g2_buf_1
X_23673_ _02046_ _03952_ VPWR VGND _03953_ sg13g2_nor2_1
X_23674_ _03814_ _03950_ _03953_ _03823_ VPWR VGND 
+ _03954_
+ sg13g2_a22oi_1
X_23675_ _03757_ VPWR VGND _03955_ sg13g2_buf_1
X_23676_ _03955_ VPWR VGND _03956_ sg13g2_buf_1
X_23677_ _03815_ VPWR VGND _03957_ sg13g2_buf_1
X_23678_ _02024_ _03827_ VPWR VGND _03958_ sg13g2_nand2b_1
X_23679_ _03957_ _02046_ _03958_ VPWR VGND _03959_ sg13g2_o21ai_1
X_23680_ _03956_ _03959_ _03831_ VPWR VGND _03960_ sg13g2_a21oi_1
X_23681_ _03948_ _03954_ _03960_ VPWR VGND _03961_ sg13g2_a21oi_1
X_23682_ _03900_ _03945_ _03947_ _03961_ VPWR VGND 
+ _03962_
+ sg13g2_nor4_1
X_23683_ _03925_ _03943_ _03962_ VPWR VGND _03963_ sg13g2_nor3_1
X_23684_ _03923_ _03963_ _03721_ VPWR VGND _03964_ sg13g2_o21ai_1
X_23685_ _03721_ _03875_ _03964_ VPWR VGND _03965_ sg13g2_o21ai_1
X_23686_ _03780_ VPWR VGND _03966_ sg13g2_buf_1
X_23687_ _03966_ VPWR VGND _03967_ sg13g2_buf_1
X_23688_ _03728_ VPWR VGND _03968_ sg13g2_buf_1
X_23689_ _03732_ VPWR VGND _03969_ sg13g2_buf_1
X_23690_ _03734_ VPWR VGND _03970_ sg13g2_buf_1
X_23691_ _03970_ VPWR VGND _03971_ sg13g2_buf_1
X_23692_ _03971_ VPWR VGND _03972_ sg13g2_buf_1
X_23693_ _02699_ VPWR VGND _03973_ sg13g2_buf_1
X_23694_ _03973_ VPWR VGND _03974_ sg13g2_buf_1
X_23695_ _03742_ VPWR VGND _03975_ sg13g2_buf_1
X_23696_ _03975_ VPWR VGND _03976_ sg13g2_buf_1
X_23697_ _02710_ VPWR VGND _03977_ sg13g2_buf_1
X_23698_ _03977_ VPWR VGND _03978_ sg13g2_buf_1
X_23699_ _03978_ _02618_ VPWR VGND _03979_ sg13g2_nor2_1
X_23700_ _02639_ _03843_ VPWR VGND _03980_ sg13g2_nor2_1
X_23701_ _02709_ VPWR VGND _03981_ sg13g2_buf_1
X_23702_ _03981_ VPWR VGND _03982_ sg13g2_buf_1
X_23703_ _03982_ VPWR VGND _03983_ sg13g2_buf_1
X_23704_ _03983_ VPWR VGND _03984_ sg13g2_buf_1
X_23705_ _03976_ _03979_ _03980_ _03984_ VPWR VGND 
+ _03985_
+ sg13g2_a22oi_1
X_23706_ _03730_ VPWR VGND _03986_ sg13g2_buf_1
X_23707_ _03986_ VPWR VGND _03987_ sg13g2_buf_1
X_23708_ _03762_ VPWR VGND _03988_ sg13g2_buf_1
X_23709_ _03988_ VPWR VGND _03989_ sg13g2_buf_1
X_23710_ _02618_ _03989_ VPWR VGND _03990_ sg13g2_nand2b_1
X_23711_ _03983_ _02639_ _03990_ VPWR VGND _03991_ sg13g2_o21ai_1
X_23712_ _03767_ VPWR VGND _03992_ sg13g2_buf_1
X_23713_ _03992_ VPWR VGND _03993_ sg13g2_buf_1
X_23714_ _03987_ _03991_ _03993_ VPWR VGND _03994_ sg13g2_a21oi_1
X_23715_ _03974_ _03985_ _03994_ VPWR VGND _03995_ sg13g2_a21oi_1
X_23716_ _00110_ _03969_ _03972_ _02660_ _03995_ VPWR 
+ VGND
+ _03996_ sg13g2_a221oi_1
X_23717_ _03774_ VPWR VGND _03997_ sg13g2_buf_1
X_23718_ \atbs_core_0.spike_memory_0.n2417_o[0]\ _03876_ VPWR VGND _03998_ sg13g2_nor2_1
X_23719_ _07563_ VPWR VGND _03999_ sg13g2_buf_1
X_23720_ _03999_ VPWR VGND _04000_ sg13g2_buf_1
X_23721_ \atbs_core_0.spike_memory_0.n2414_o[0]\ _04000_ _03722_ VPWR VGND _04001_ sg13g2_o21ai_1
X_23722_ _02699_ VPWR VGND _04002_ sg13g2_buf_1
X_23723_ _03742_ VPWR VGND _04003_ sg13g2_buf_1
X_23724_ _02710_ VPWR VGND _04004_ sg13g2_buf_1
X_23725_ _04004_ _12572_ VPWR VGND _04005_ sg13g2_nor2_1
X_23726_ _03749_ VPWR VGND _04006_ sg13g2_buf_1
X_23727_ _12595_ _04006_ VPWR VGND _04007_ sg13g2_nor2_1
X_23728_ _04003_ _04005_ _04007_ _03978_ VPWR VGND 
+ _04008_
+ sg13g2_a22oi_1
X_23729_ _03730_ VPWR VGND _04009_ sg13g2_buf_1
X_23730_ _04009_ VPWR VGND _04010_ sg13g2_buf_1
X_23731_ _03762_ VPWR VGND _04011_ sg13g2_buf_1
X_23732_ _12572_ _04011_ VPWR VGND _04012_ sg13g2_nand2b_1
X_23733_ _03977_ _12595_ _04012_ VPWR VGND _04013_ sg13g2_o21ai_1
X_23734_ _04010_ _04013_ _03839_ VPWR VGND _04014_ sg13g2_a21oi_1
X_23735_ _04002_ _04008_ _04014_ VPWR VGND _04015_ sg13g2_a21oi_1
X_23736_ _03998_ _04001_ _04015_ VPWR VGND _04016_ sg13g2_or3_1
X_23737_ _03997_ _04016_ VPWR VGND _04017_ sg13g2_nand2_1
X_23738_ _03968_ _03996_ _04017_ VPWR VGND _04018_ sg13g2_o21ai_1
X_23739_ \atbs_core_0.spike_memory_0.n2413_o[0]\ _12087_ VPWR VGND _04019_ sg13g2_nor2_1
X_23740_ \atbs_core_0.spike_memory_0.n2410_o[0]\ _03836_ VPWR VGND _04020_ sg13g2_nor2_1
X_23741_ _02700_ VPWR VGND _04021_ sg13g2_buf_1
X_23742_ _03882_ _12516_ VPWR VGND _04022_ sg13g2_nor2_1
X_23743_ _03785_ VPWR VGND _04023_ sg13g2_buf_1
X_23744_ _12540_ _04023_ VPWR VGND _04024_ sg13g2_nor2_1
X_23745_ _03881_ _04022_ _04024_ _03887_ VPWR VGND 
+ _04025_
+ sg13g2_a22oi_1
X_23746_ _03791_ VPWR VGND _04026_ sg13g2_buf_1
X_23747_ _12516_ _04026_ VPWR VGND _04027_ sg13g2_nand2b_1
X_23748_ _03886_ _12540_ _04027_ VPWR VGND _04028_ sg13g2_o21ai_1
X_23749_ _03759_ _04028_ _03895_ VPWR VGND _04029_ sg13g2_a21oi_1
X_23750_ _04021_ _04025_ _04029_ VPWR VGND _04030_ sg13g2_a21oi_1
X_23751_ _04019_ _04020_ _04030_ VPWR VGND _04031_ sg13g2_nor3_1
X_23752_ _03779_ VPWR VGND _04032_ sg13g2_buf_1
X_23753_ \atbs_core_0.spike_memory_0.n2436_q[1197]\ _03971_ VPWR VGND _04033_ sg13g2_nand2b_1
X_23754_ \atbs_core_0.spike_memory_0.n2418_o[0]\ _04032_ _04033_ VPWR VGND _04034_ sg13g2_o21ai_1
X_23755_ _03813_ VPWR VGND _04035_ sg13g2_buf_1
X_23756_ _03816_ _12627_ VPWR VGND _04036_ sg13g2_nor2_1
X_23757_ _12653_ _03819_ VPWR VGND _04037_ sg13g2_nor2_1
X_23758_ _04035_ _04036_ _04037_ _03823_ VPWR VGND 
+ _04038_
+ sg13g2_a22oi_1
X_23759_ _12627_ _03916_ VPWR VGND _04039_ sg13g2_nand2b_1
X_23760_ _03930_ _12653_ _04039_ VPWR VGND _04040_ sg13g2_o21ai_1
X_23761_ _03825_ _04040_ _03831_ VPWR VGND _04041_ sg13g2_a21oi_1
X_23762_ _03905_ _04038_ _04041_ VPWR VGND _04042_ sg13g2_a21oi_1
X_23763_ _04034_ _04042_ _03997_ VPWR VGND _04043_ sg13g2_o21ai_1
X_23764_ _03801_ _04031_ _04043_ VPWR VGND _04044_ sg13g2_o21ai_1
X_23765_ _03720_ VPWR VGND _04045_ sg13g2_buf_1
X_23766_ _03967_ _04018_ _04044_ _04016_ _04045_ VPWR 
+ VGND
+ _04046_ sg13g2_a221oi_1
X_23767_ _03842_ VPWR VGND _04047_ sg13g2_buf_1
X_23768_ _03855_ _02134_ VPWR VGND _04048_ sg13g2_nor2_1
X_23769_ _02157_ _03951_ VPWR VGND _04049_ sg13g2_nor2_1
X_23770_ _03845_ VPWR VGND _04050_ sg13g2_buf_1
X_23771_ _04050_ VPWR VGND _04051_ sg13g2_buf_1
X_23772_ _04051_ VPWR VGND _04052_ sg13g2_buf_1
X_23773_ _04047_ _04048_ _04049_ _04052_ VPWR VGND 
+ _04053_
+ sg13g2_a22oi_1
X_23774_ _03862_ VPWR VGND _04054_ sg13g2_buf_1
X_23775_ _02134_ _04054_ VPWR VGND _04055_ sg13g2_nand2b_1
X_23776_ _03815_ _02157_ _04055_ VPWR VGND _04056_ sg13g2_o21ai_1
X_23777_ _03955_ _04056_ _03868_ VPWR VGND _04057_ sg13g2_a21oi_1
X_23778_ _03993_ _04053_ _04057_ VPWR VGND _04058_ sg13g2_a21oi_1
X_23779_ _00112_ _03732_ _03736_ _02180_ _04058_ VPWR 
+ VGND
+ _04059_ sg13g2_a221oi_1
X_23780_ \atbs_core_0.spike_memory_0.n2385_o[0]\ _03802_ VPWR VGND _04060_ sg13g2_nor2_1
X_23781_ \atbs_core_0.spike_memory_0.n2382_o[0]\ _03778_ _07552_ VPWR VGND _04061_ sg13g2_o21ai_1
X_23782_ _03749_ VPWR VGND _04062_ sg13g2_buf_1
X_23783_ _03846_ _02286_ VPWR VGND _04063_ sg13g2_nor2_1
X_23784_ _02309_ _03850_ VPWR VGND _04064_ sg13g2_nor2_1
X_23785_ _04062_ _04063_ _04064_ _03855_ VPWR VGND 
+ _04065_
+ sg13g2_a22oi_1
X_23786_ _02286_ _03862_ VPWR VGND _04066_ sg13g2_nand2b_1
X_23787_ _03854_ _02309_ _04066_ VPWR VGND _04067_ sg13g2_o21ai_1
X_23788_ _02698_ VPWR VGND _04068_ sg13g2_buf_1
X_23789_ _03859_ _04067_ _04068_ VPWR VGND _04069_ sg13g2_a21oi_1
X_23790_ _03839_ _04065_ _04069_ VPWR VGND _04070_ sg13g2_a21oi_1
X_23791_ _04060_ _04061_ _04070_ VPWR VGND _04071_ sg13g2_or3_1
X_23792_ _03774_ _04071_ VPWR VGND _04072_ sg13g2_nand2_1
X_23793_ _03926_ _04059_ _04072_ VPWR VGND _04073_ sg13g2_o21ai_1
X_23794_ _03800_ VPWR VGND _04074_ sg13g2_buf_1
X_23795_ _12084_ VPWR VGND _04075_ sg13g2_buf_1
X_23796_ _04075_ VPWR VGND _04076_ sg13g2_buf_1
X_23797_ \atbs_core_0.spike_memory_0.n2381_o[0]\ _04076_ VPWR VGND _04077_ sg13g2_nor2_1
X_23798_ _07563_ VPWR VGND _04078_ sg13g2_buf_1
X_23799_ _04078_ VPWR VGND _04079_ sg13g2_buf_1
X_23800_ \atbs_core_0.spike_memory_0.n2378_o[0]\ _04079_ VPWR VGND _04080_ sg13g2_nor2_1
X_23801_ _03768_ VPWR VGND _04081_ sg13g2_buf_1
X_23802_ _03785_ VPWR VGND _04082_ sg13g2_buf_1
X_23803_ _04011_ VPWR VGND _04083_ sg13g2_buf_1
X_23804_ _04083_ _02231_ VPWR VGND _04084_ sg13g2_nor2_1
X_23805_ _03741_ VPWR VGND _04085_ sg13g2_buf_1
X_23806_ _04085_ VPWR VGND _04086_ sg13g2_buf_1
X_23807_ _02254_ _04086_ VPWR VGND _04087_ sg13g2_nor2_1
X_23808_ _03762_ VPWR VGND _04088_ sg13g2_buf_1
X_23809_ _04088_ VPWR VGND _04089_ sg13g2_buf_1
X_23810_ _04089_ VPWR VGND _04090_ sg13g2_buf_1
X_23811_ _04082_ _04084_ _04087_ _04090_ VPWR VGND 
+ _04091_
+ sg13g2_a22oi_1
X_23812_ _03859_ VPWR VGND _04092_ sg13g2_buf_1
X_23813_ _02709_ VPWR VGND _04093_ sg13g2_buf_1
X_23814_ _04093_ VPWR VGND _04094_ sg13g2_buf_1
X_23815_ _02231_ _04094_ VPWR VGND _04095_ sg13g2_nand2b_1
X_23816_ _04089_ _02254_ _04095_ VPWR VGND _04096_ sg13g2_o21ai_1
X_23817_ _02698_ VPWR VGND _04097_ sg13g2_buf_1
X_23818_ _04097_ VPWR VGND _04098_ sg13g2_buf_1
X_23819_ _04092_ _04096_ _04098_ VPWR VGND _04099_ sg13g2_a21oi_1
X_23820_ _04081_ _04091_ _04099_ VPWR VGND _04100_ sg13g2_a21oi_1
X_23821_ _04077_ _04080_ _04100_ VPWR VGND _04101_ sg13g2_nor3_1
X_23822_ _04078_ VPWR VGND _04102_ sg13g2_buf_1
X_23823_ \atbs_core_0.spike_memory_0.n2389_o[0]\ _03735_ VPWR VGND _04103_ sg13g2_nand2b_1
X_23824_ \atbs_core_0.spike_memory_0.n2386_o[0]\ _04102_ _04103_ VPWR VGND _04104_ sg13g2_o21ai_1
X_23825_ _03763_ VPWR VGND _04105_ sg13g2_buf_1
X_23826_ _04105_ _02342_ VPWR VGND _04106_ sg13g2_nor2_1
X_23827_ _03741_ VPWR VGND _04107_ sg13g2_buf_1
X_23828_ _04107_ VPWR VGND _04108_ sg13g2_buf_1
X_23829_ _02366_ _04108_ VPWR VGND _04109_ sg13g2_nor2_1
X_23830_ _03762_ VPWR VGND _04110_ sg13g2_buf_1
X_23831_ _04110_ VPWR VGND _04111_ sg13g2_buf_1
X_23832_ _04111_ VPWR VGND _04112_ sg13g2_buf_1
X_23833_ _03932_ _04106_ _04109_ _04112_ VPWR VGND 
+ _04113_
+ sg13g2_a22oi_1
X_23834_ _03986_ VPWR VGND _04114_ sg13g2_buf_1
X_23835_ _03745_ VPWR VGND _04115_ sg13g2_buf_1
X_23836_ _02342_ _04115_ VPWR VGND _04116_ sg13g2_nand2b_1
X_23837_ _03764_ _02366_ _04116_ VPWR VGND _04117_ sg13g2_o21ai_1
X_23838_ _02699_ VPWR VGND _04118_ sg13g2_buf_1
X_23839_ _04114_ _04117_ _04118_ VPWR VGND _04119_ sg13g2_a21oi_1
X_23840_ _03919_ _04113_ _04119_ VPWR VGND _04120_ sg13g2_a21oi_1
X_23841_ _04104_ _04120_ _03728_ VPWR VGND _04121_ sg13g2_o21ai_1
X_23842_ _04074_ _04101_ _04121_ VPWR VGND _04122_ sg13g2_o21ai_1
X_23843_ _03967_ _04073_ _04122_ _04071_ VPWR VGND 
+ _04123_
+ sg13g2_a22oi_1
X_23844_ _04045_ _04123_ VPWR VGND _04124_ sg13g2_and2_1
X_23845_ _03718_ _04046_ _04124_ VPWR VGND _04125_ sg13g2_nor3_1
X_23846_ _03719_ _03965_ _04125_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[0]\ sg13g2_a21oi_1
X_23847_ _03900_ VPWR VGND _04126_ sg13g2_buf_1
X_23848_ _03882_ _02401_ VPWR VGND _04127_ sg13g2_nor2_1
X_23849_ _02420_ _04023_ VPWR VGND _04128_ sg13g2_nor2_1
X_23850_ _03881_ _04127_ _04128_ _03887_ VPWR VGND 
+ _04129_
+ sg13g2_a22oi_1
X_23851_ _02401_ _04026_ VPWR VGND _04130_ sg13g2_nand2b_1
X_23852_ _03886_ _02420_ _04130_ VPWR VGND _04131_ sg13g2_o21ai_1
X_23853_ _03889_ _04131_ _03895_ VPWR VGND _04132_ sg13g2_a21oi_1
X_23854_ _03880_ _04129_ _04132_ VPWR VGND _04133_ sg13g2_a21oi_1
X_23855_ _00141_ _03733_ _03737_ _02452_ _04133_ VPWR 
+ VGND
+ _04134_ sg13g2_a221oi_1
X_23856_ \atbs_core_0.spike_memory_0.n2401_o[10]\ _03901_ VPWR VGND _04135_ sg13g2_nor2_1
X_23857_ \atbs_core_0.spike_memory_0.n2398_o[10]\ _03903_ VPWR VGND _04136_ sg13g2_nor2_1
X_23858_ _03907_ _02534_ VPWR VGND _04137_ sg13g2_nor2_1
X_23859_ _02555_ _03909_ VPWR VGND _04138_ sg13g2_nor2_1
X_23860_ _03906_ _04137_ _04138_ _03911_ VPWR VGND 
+ _04139_
+ sg13g2_a22oi_1
X_23861_ _02534_ _03916_ VPWR VGND _04140_ sg13g2_nand2b_1
X_23862_ _03930_ _02555_ _04140_ VPWR VGND _04141_ sg13g2_o21ai_1
X_23863_ _03830_ VPWR VGND _04142_ sg13g2_buf_1
X_23864_ _03913_ _04141_ _04142_ VPWR VGND _04143_ sg13g2_a21oi_1
X_23865_ _03905_ _04139_ _04143_ VPWR VGND _04144_ sg13g2_a21oi_1
X_23866_ _03900_ _04135_ _04136_ _04144_ VPWR VGND 
+ _04145_
+ sg13g2_nor4_1
X_23867_ _04126_ _04134_ _04145_ VPWR VGND _04146_ sg13g2_a21oi_1
X_23868_ \atbs_core_0.spike_memory_0.n2397_o[10]\ _12087_ VPWR VGND _04147_ sg13g2_nor2_1
X_23869_ \atbs_core_0.spike_memory_0.n2394_o[10]\ _03903_ VPWR VGND _04148_ sg13g2_nor2_1
X_23870_ _02700_ VPWR VGND _04149_ sg13g2_buf_1
X_23871_ _03813_ VPWR VGND _04150_ sg13g2_buf_1
X_23872_ _03826_ _02487_ VPWR VGND _04151_ sg13g2_nor2_1
X_23873_ _03818_ VPWR VGND _04152_ sg13g2_buf_1
X_23874_ _02508_ _04152_ VPWR VGND _04153_ sg13g2_nor2_1
X_23875_ _03914_ VPWR VGND _04154_ sg13g2_buf_1
X_23876_ _04150_ _04151_ _04153_ _04154_ VPWR VGND 
+ _04155_
+ sg13g2_a22oi_1
X_23877_ _02487_ _03937_ VPWR VGND _04156_ sg13g2_nand2b_1
X_23878_ _02712_ _02508_ _04156_ VPWR VGND _04157_ sg13g2_o21ai_1
X_23879_ _03830_ VPWR VGND _04158_ sg13g2_buf_1
X_23880_ _03936_ _04157_ _04158_ VPWR VGND _04159_ sg13g2_a21oi_1
X_23881_ _04149_ _04155_ _04159_ VPWR VGND _04160_ sg13g2_a21oi_1
X_23882_ _03926_ _04147_ _04148_ _04160_ VPWR VGND 
+ _04161_
+ sg13g2_nor4_1
X_23883_ \atbs_core_0.spike_memory_0.n2405_o[10]\ _03944_ VPWR VGND _04162_ sg13g2_nor2_1
X_23884_ \atbs_core_0.spike_memory_0.n2402_o[10]\ _03946_ VPWR VGND _04163_ sg13g2_nor2_1
X_23885_ _03949_ _02582_ VPWR VGND _04164_ sg13g2_nor2_1
X_23886_ _02603_ _03952_ VPWR VGND _04165_ sg13g2_nor2_1
X_23887_ _03814_ _04164_ _04165_ _03823_ VPWR VGND 
+ _04166_
+ sg13g2_a22oi_1
X_23888_ _03915_ VPWR VGND _04167_ sg13g2_buf_1
X_23889_ _02582_ _04167_ VPWR VGND _04168_ sg13g2_nand2b_1
X_23890_ _03957_ _02603_ _04168_ VPWR VGND _04169_ sg13g2_o21ai_1
X_23891_ _03956_ _04169_ _03831_ VPWR VGND _04170_ sg13g2_a21oi_1
X_23892_ _03948_ _04166_ _04170_ VPWR VGND _04171_ sg13g2_a21oi_1
X_23893_ _03900_ _04162_ _04163_ _04171_ VPWR VGND 
+ _04172_
+ sg13g2_nor4_1
X_23894_ _03967_ _04161_ _04172_ VPWR VGND _04173_ sg13g2_nor3_1
X_23895_ _03725_ _04146_ _04173_ VPWR VGND _04174_ sg13g2_a21oi_1
X_23896_ \atbs_core_0.spike_memory_0.n2365_o[10]\ _03877_ VPWR VGND _04175_ sg13g2_nor2_1
X_23897_ \atbs_core_0.spike_memory_0.n2362_o[10]\ _03836_ VPWR VGND _04176_ sg13g2_nor2_1
X_23898_ _03882_ _12565_ VPWR VGND _04177_ sg13g2_nor2_1
X_23899_ _02010_ _04023_ VPWR VGND _04178_ sg13g2_nor2_1
X_23900_ _03881_ _04177_ _04178_ _03887_ VPWR VGND 
+ _04179_
+ sg13g2_a22oi_1
X_23901_ _12565_ _04026_ VPWR VGND _04180_ sg13g2_nand2b_1
X_23902_ _03886_ _02010_ _04180_ VPWR VGND _04181_ sg13g2_o21ai_1
X_23903_ _03889_ _04181_ _03895_ VPWR VGND _04182_ sg13g2_a21oi_1
X_23904_ _03880_ _04179_ _04182_ VPWR VGND _04183_ sg13g2_a21oi_1
X_23905_ _03728_ _04175_ _04176_ _04183_ VPWR VGND 
+ _04184_
+ sg13g2_nor4_1
X_23906_ \atbs_core_0.spike_memory_0.n2373_o[10]\ _03901_ VPWR VGND _04185_ sg13g2_nor2_1
X_23907_ \atbs_core_0.spike_memory_0.n2370_o[10]\ _03903_ VPWR VGND _04186_ sg13g2_nor2_1
X_23908_ _03907_ _02091_ VPWR VGND _04187_ sg13g2_nor2_1
X_23909_ _02114_ _03909_ VPWR VGND _04188_ sg13g2_nor2_1
X_23910_ _03906_ _04187_ _04188_ _03911_ VPWR VGND 
+ _04189_
+ sg13g2_a22oi_1
X_23911_ _02091_ _03916_ VPWR VGND _04190_ sg13g2_nand2b_1
X_23912_ _03914_ _02114_ _04190_ VPWR VGND _04191_ sg13g2_o21ai_1
X_23913_ _03913_ _04191_ _03919_ VPWR VGND _04192_ sg13g2_a21oi_1
X_23914_ _03905_ _04189_ _04192_ VPWR VGND _04193_ sg13g2_a21oi_1
X_23915_ _03900_ _04185_ _04186_ _04193_ VPWR VGND 
+ _04194_
+ sg13g2_nor4_1
X_23916_ _03724_ _04184_ _04194_ VPWR VGND _04195_ sg13g2_nor3_1
X_23917_ \atbs_core_0.spike_memory_0.n2361_o[10]\ _12087_ VPWR VGND _04196_ sg13g2_nor2_1
X_23918_ \atbs_core_0.spike_memory_0.n2358_o[10]\ _03903_ VPWR VGND _04197_ sg13g2_nor2_1
X_23919_ _03930_ _02129_ VPWR VGND _04198_ sg13g2_nor2_1
X_23920_ _02304_ _03932_ VPWR VGND _04199_ sg13g2_nor2_1
X_23921_ _03929_ _04198_ _04199_ _02713_ VPWR VGND 
+ _04200_
+ sg13g2_a22oi_1
X_23922_ _02129_ _03937_ VPWR VGND _04201_ sg13g2_nand2b_1
X_23923_ _02712_ _02304_ _04201_ VPWR VGND _04202_ sg13g2_o21ai_1
X_23924_ _03936_ _04202_ _03940_ VPWR VGND _04203_ sg13g2_a21oi_1
X_23925_ _02701_ _04200_ _04203_ VPWR VGND _04204_ sg13g2_a21oi_1
X_23926_ _03728_ _04196_ _04197_ _04204_ VPWR VGND 
+ _04205_
+ sg13g2_nor4_1
X_23927_ \atbs_core_0.spike_memory_0.n2369_o[10]\ _03901_ VPWR VGND _04206_ sg13g2_nor2_1
X_23928_ \atbs_core_0.spike_memory_0.n2366_o[10]\ _03807_ VPWR VGND _04207_ sg13g2_nor2_1
X_23929_ _03949_ _02036_ VPWR VGND _04208_ sg13g2_nor2_1
X_23930_ _02059_ _03952_ VPWR VGND _04209_ sg13g2_nor2_1
X_23931_ _03814_ _04208_ _04209_ _03823_ VPWR VGND 
+ _04210_
+ sg13g2_a22oi_1
X_23932_ _02036_ _03827_ VPWR VGND _04211_ sg13g2_nand2b_1
X_23933_ _03957_ _02059_ _04211_ VPWR VGND _04212_ sg13g2_o21ai_1
X_23934_ _03825_ _04212_ _03831_ VPWR VGND _04213_ sg13g2_a21oi_1
X_23935_ _03948_ _04210_ _04213_ VPWR VGND _04214_ sg13g2_a21oi_1
X_23936_ _03900_ _04206_ _04207_ _04214_ VPWR VGND 
+ _04215_
+ sg13g2_nor4_1
X_23937_ _03925_ _04205_ _04215_ VPWR VGND _04216_ sg13g2_nor3_1
X_23938_ _04195_ _04216_ _03721_ VPWR VGND _04217_ sg13g2_o21ai_1
X_23939_ _03721_ _04174_ _04217_ VPWR VGND _04218_ sg13g2_o21ai_1
X_23940_ _03899_ VPWR VGND _04219_ sg13g2_buf_1
X_23941_ _04083_ _02629_ VPWR VGND _04220_ sg13g2_nor2_1
X_23942_ _02650_ _04086_ VPWR VGND _04221_ sg13g2_nor2_1
X_23943_ _04082_ _04220_ _04221_ _04090_ VPWR VGND 
+ _04222_
+ sg13g2_a22oi_1
X_23944_ _02629_ _04094_ VPWR VGND _04223_ sg13g2_nand2b_1
X_23945_ _04089_ _02650_ _04223_ VPWR VGND _04224_ sg13g2_o21ai_1
X_23946_ _04092_ _04224_ _04098_ VPWR VGND _04225_ sg13g2_a21oi_1
X_23947_ _04081_ _04222_ _04225_ VPWR VGND _04226_ sg13g2_a21oi_1
X_23948_ _00140_ _03732_ _03736_ _02680_ _04226_ VPWR 
+ VGND
+ _04227_ sg13g2_a221oi_1
X_23949_ \atbs_core_0.spike_memory_0.n2417_o[10]\ _04076_ VPWR VGND _04228_ sg13g2_nor2_1
X_23950_ _03999_ VPWR VGND _04229_ sg13g2_buf_1
X_23951_ _04229_ VPWR VGND _04230_ sg13g2_buf_1
X_23952_ \atbs_core_0.spike_memory_0.n2414_o[10]\ _04230_ VPWR VGND _04231_ sg13g2_nor2_1
X_23953_ _04105_ _12584_ VPWR VGND _04232_ sg13g2_nor2_1
X_23954_ _12607_ _04108_ VPWR VGND _04233_ sg13g2_nor2_1
X_23955_ _03932_ _04232_ _04233_ _04112_ VPWR VGND 
+ _04234_
+ sg13g2_a22oi_1
X_23956_ _03986_ VPWR VGND _04235_ sg13g2_buf_1
X_23957_ _03763_ VPWR VGND _04236_ sg13g2_buf_1
X_23958_ _02710_ VPWR VGND _04237_ sg13g2_buf_1
X_23959_ _12584_ _04237_ VPWR VGND _04238_ sg13g2_nand2b_1
X_23960_ _04236_ _12607_ _04238_ VPWR VGND _04239_ sg13g2_o21ai_1
X_23961_ _04235_ _04239_ _03973_ VPWR VGND _04240_ sg13g2_a21oi_1
X_23962_ _04158_ _04234_ _04240_ VPWR VGND _04241_ sg13g2_a21oi_1
X_23963_ _03899_ _04228_ _04231_ _04241_ VPWR VGND 
+ _04242_
+ sg13g2_nor4_1
X_23964_ _04219_ _04227_ _04242_ VPWR VGND _04243_ sg13g2_a21oi_1
X_23965_ _03773_ VPWR VGND _04244_ sg13g2_buf_1
X_23966_ _03802_ VPWR VGND _04245_ sg13g2_buf_1
X_23967_ \atbs_core_0.spike_memory_0.n2413_o[10]\ _04245_ VPWR VGND _04246_ sg13g2_nor2_1
X_23968_ _04078_ VPWR VGND _04247_ sg13g2_buf_1
X_23969_ \atbs_core_0.spike_memory_0.n2410_o[10]\ _04247_ VPWR VGND _04248_ sg13g2_nor2_1
X_23970_ _04083_ _12529_ VPWR VGND _04249_ sg13g2_nor2_1
X_23971_ _04107_ VPWR VGND _04250_ sg13g2_buf_1
X_23972_ _12552_ _04250_ VPWR VGND _04251_ sg13g2_nor2_1
X_23973_ _04023_ _04249_ _04251_ _04090_ VPWR VGND 
+ _04252_
+ sg13g2_a22oi_1
X_23974_ _03986_ VPWR VGND _04253_ sg13g2_buf_1
X_23975_ _04093_ VPWR VGND _04254_ sg13g2_buf_1
X_23976_ _12529_ _04254_ VPWR VGND _04255_ sg13g2_nand2b_1
X_23977_ _04089_ _12552_ _04255_ VPWR VGND _04256_ sg13g2_o21ai_1
X_23978_ _04253_ _04256_ _04098_ VPWR VGND _04257_ sg13g2_a21oi_1
X_23979_ _04081_ _04252_ _04257_ VPWR VGND _04258_ sg13g2_a21oi_1
X_23980_ _04244_ _04246_ _04248_ _04258_ VPWR VGND 
+ _04259_
+ sg13g2_nor4_1
X_23981_ _04075_ VPWR VGND _04260_ sg13g2_buf_1
X_23982_ \atbs_core_0.spike_memory_0.n2436_q[1207]\ _04260_ VPWR VGND _04261_ sg13g2_nor2_1
X_23983_ \atbs_core_0.spike_memory_0.n2418_o[10]\ _04079_ VPWR VGND _04262_ sg13g2_nor2_1
X_23984_ _03768_ VPWR VGND _04263_ sg13g2_buf_1
X_23985_ _04111_ _12641_ VPWR VGND _04264_ sg13g2_nor2_1
X_23986_ _04107_ VPWR VGND _04265_ sg13g2_buf_1
X_23987_ _12666_ _04265_ VPWR VGND _04266_ sg13g2_nor2_1
X_23988_ _04011_ VPWR VGND _04267_ sg13g2_buf_1
X_23989_ _04267_ VPWR VGND _04268_ sg13g2_buf_1
X_23990_ _03884_ _04264_ _04266_ _04268_ VPWR VGND 
+ _04269_
+ sg13g2_a22oi_1
X_23991_ _12641_ _04004_ VPWR VGND _04270_ sg13g2_nand2b_1
X_23992_ _04267_ _12666_ _04270_ VPWR VGND _04271_ sg13g2_o21ai_1
X_23993_ _02699_ VPWR VGND _04272_ sg13g2_buf_1
X_23994_ _04235_ _04271_ _04272_ VPWR VGND _04273_ sg13g2_a21oi_1
X_23995_ _04263_ _04269_ _04273_ VPWR VGND _04274_ sg13g2_a21oi_1
X_23996_ _03899_ _04261_ _04262_ _04274_ VPWR VGND 
+ _04275_
+ sg13g2_nor4_1
X_23997_ _12090_ VPWR VGND _04276_ sg13g2_buf_1
X_23998_ _04276_ VPWR VGND _04277_ sg13g2_buf_1
X_23999_ _04259_ _04275_ _04277_ VPWR VGND _04278_ sg13g2_o21ai_1
X_24000_ _03925_ _04243_ _04278_ VPWR VGND _04279_ sg13g2_o21ai_1
X_24001_ _04006_ VPWR VGND _04280_ sg13g2_buf_1
X_24002_ _03989_ _02146_ VPWR VGND _04281_ sg13g2_nor2_1
X_24003_ _02169_ _03851_ VPWR VGND _04282_ sg13g2_nor2_1
X_24004_ _03847_ VPWR VGND _04283_ sg13g2_buf_1
X_24005_ _04280_ _04281_ _04282_ _04283_ VPWR VGND 
+ _04284_
+ sg13g2_a22oi_1
X_24006_ _02146_ _03982_ VPWR VGND _04285_ sg13g2_nand2b_1
X_24007_ _03847_ _02169_ _04285_ VPWR VGND _04286_ sg13g2_o21ai_1
X_24008_ _04068_ VPWR VGND _04287_ sg13g2_buf_1
X_24009_ _03860_ _04286_ _04287_ VPWR VGND _04288_ sg13g2_a21oi_1
X_24010_ _03840_ _04284_ _04288_ VPWR VGND _04289_ sg13g2_a21oi_1
X_24011_ _00142_ _03732_ _03736_ _02207_ _04289_ VPWR 
+ VGND
+ _04290_ sg13g2_a221oi_1
X_24012_ \atbs_core_0.spike_memory_0.n2385_o[10]\ _03802_ VPWR VGND _04291_ sg13g2_nor2_1
X_24013_ _07563_ VPWR VGND _04292_ sg13g2_buf_1
X_24014_ \atbs_core_0.spike_memory_0.n2382_o[10]\ _04292_ _07552_ VPWR VGND _04293_ sg13g2_o21ai_1
X_24015_ _03767_ VPWR VGND _04294_ sg13g2_buf_1
X_24016_ _04011_ _02298_ VPWR VGND _04295_ sg13g2_nor2_1
X_24017_ _02321_ _04085_ VPWR VGND _04296_ sg13g2_nor2_1
X_24018_ _03750_ _04295_ _04296_ _03989_ VPWR VGND 
+ _04297_
+ sg13g2_a22oi_1
X_24019_ _02298_ _04093_ VPWR VGND _04298_ sg13g2_nand2b_1
X_24020_ _03988_ _02321_ _04298_ VPWR VGND _04299_ sg13g2_o21ai_1
X_24021_ _03859_ _04299_ _04097_ VPWR VGND _04300_ sg13g2_a21oi_1
X_24022_ _04294_ _04297_ _04300_ VPWR VGND _04301_ sg13g2_a21oi_1
X_24023_ _04291_ _04293_ _04301_ VPWR VGND _04302_ sg13g2_or3_1
X_24024_ _03728_ _04302_ VPWR VGND _04303_ sg13g2_nand2_1
X_24025_ _03926_ _04290_ _04303_ VPWR VGND _04304_ sg13g2_o21ai_1
X_24026_ \atbs_core_0.spike_memory_0.n2381_o[10]\ _04076_ VPWR VGND _04305_ sg13g2_nor2_1
X_24027_ \atbs_core_0.spike_memory_0.n2378_o[10]\ _04230_ VPWR VGND _04306_ sg13g2_nor2_1
X_24028_ _04105_ _02243_ VPWR VGND _04307_ sg13g2_nor2_1
X_24029_ _02266_ _04108_ VPWR VGND _04308_ sg13g2_nor2_1
X_24030_ _03932_ _04307_ _04308_ _04112_ VPWR VGND 
+ _04309_
+ sg13g2_a22oi_1
X_24031_ _02243_ _04237_ VPWR VGND _04310_ sg13g2_nand2b_1
X_24032_ _04111_ _02266_ _04310_ VPWR VGND _04311_ sg13g2_o21ai_1
X_24033_ _04114_ _04311_ _03973_ VPWR VGND _04312_ sg13g2_a21oi_1
X_24034_ _04158_ _04309_ _04312_ VPWR VGND _04313_ sg13g2_a21oi_1
X_24035_ _04305_ _04306_ _04313_ VPWR VGND _04314_ sg13g2_nor3_1
X_24036_ \atbs_core_0.spike_memory_0.n2389_o[10]\ _03735_ VPWR VGND _04315_ sg13g2_nand2b_1
X_24037_ \atbs_core_0.spike_memory_0.n2386_o[10]\ _04247_ _04315_ VPWR VGND _04316_ sg13g2_o21ai_1
X_24038_ _03868_ VPWR VGND _04317_ sg13g2_buf_1
X_24039_ _03937_ _02354_ VPWR VGND _04318_ sg13g2_nor2_1
X_24040_ _02377_ _04003_ VPWR VGND _04319_ sg13g2_nor2_1
X_24041_ _03892_ VPWR VGND _04320_ sg13g2_buf_1
X_24042_ _03952_ _04318_ _04319_ _04320_ VPWR VGND 
+ _04321_
+ sg13g2_a22oi_1
X_24043_ _02354_ _02711_ VPWR VGND _04322_ sg13g2_nand2b_1
X_24044_ _03892_ _02377_ _04322_ VPWR VGND _04323_ sg13g2_o21ai_1
X_24045_ _03738_ VPWR VGND _04324_ sg13g2_buf_1
X_24046_ _04114_ _04323_ _04324_ VPWR VGND _04325_ sg13g2_a21oi_1
X_24047_ _04317_ _04321_ _04325_ VPWR VGND _04326_ sg13g2_a21oi_1
X_24048_ _04316_ _04326_ _03728_ VPWR VGND _04327_ sg13g2_o21ai_1
X_24049_ _04074_ _04314_ _04327_ VPWR VGND _04328_ sg13g2_o21ai_1
X_24050_ _03967_ _04304_ _04328_ _04302_ VPWR VGND 
+ _04329_
+ sg13g2_a22oi_1
X_24051_ _03720_ VPWR VGND _04330_ sg13g2_buf_1
X_24052_ _04279_ _04329_ _04330_ VPWR VGND _04331_ sg13g2_mux2_1
X_24053_ _03719_ _04331_ VPWR VGND _04332_ sg13g2_nor2_1
X_24054_ _03719_ _04218_ _04332_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[10]\ sg13g2_a21oi_1
X_24055_ _07549_ VPWR VGND _04333_ sg13g2_buf_1
X_24056_ _12090_ _03727_ VPWR VGND _04334_ sg13g2_nor2_1
X_24057_ _04334_ VPWR VGND _04335_ sg13g2_buf_1
X_24058_ _04335_ VPWR VGND _04336_ sg13g2_buf_1
X_24059_ _03717_ VPWR VGND _04337_ sg13g2_buf_1
X_24060_ _03940_ VPWR VGND _04338_ sg13g2_buf_1
X_24061_ _03819_ VPWR VGND _04339_ sg13g2_buf_1
X_24062_ _03892_ VPWR VGND _04340_ sg13g2_buf_1
X_24063_ _04340_ _02402_ VPWR VGND _04341_ sg13g2_nor2_1
X_24064_ _02421_ _03976_ VPWR VGND _04342_ sg13g2_nor2_1
X_24065_ _04283_ VPWR VGND _04343_ sg13g2_buf_1
X_24066_ _04339_ _04341_ _04342_ _04343_ VPWR VGND 
+ _04344_
+ sg13g2_a22oi_1
X_24067_ _04114_ VPWR VGND _04345_ sg13g2_buf_1
X_24068_ _03763_ VPWR VGND _04346_ sg13g2_buf_1
X_24069_ _04346_ VPWR VGND _04347_ sg13g2_buf_1
X_24070_ _02402_ _03788_ VPWR VGND _04348_ sg13g2_nand2b_1
X_24071_ _04347_ _02421_ _04348_ VPWR VGND _04349_ sg13g2_o21ai_1
X_24072_ _04345_ _04349_ _03974_ VPWR VGND _04350_ sg13g2_a21oi_1
X_24073_ _04338_ _04344_ _04350_ VPWR VGND _04351_ sg13g2_a21oi_1
X_24074_ _00144_ _03733_ _03737_ _02454_ _04351_ VPWR 
+ VGND
+ _04352_ sg13g2_a221oi_1
X_24075_ _03732_ VPWR VGND _04353_ sg13g2_buf_1
X_24076_ _03972_ VPWR VGND _04354_ sg13g2_buf_1
X_24077_ _04317_ VPWR VGND _04355_ sg13g2_buf_1
X_24078_ _03952_ VPWR VGND _04356_ sg13g2_buf_1
X_24079_ _03827_ VPWR VGND _04357_ sg13g2_buf_1
X_24080_ _04357_ _02147_ VPWR VGND _04358_ sg13g2_nor2_1
X_24081_ _03782_ VPWR VGND _04359_ sg13g2_buf_1
X_24082_ _02171_ _04359_ VPWR VGND _04360_ sg13g2_nor2_1
X_24083_ _03892_ VPWR VGND _04361_ sg13g2_buf_1
X_24084_ _04361_ VPWR VGND _04362_ sg13g2_buf_1
X_24085_ _04356_ _04358_ _04360_ _04362_ VPWR VGND 
+ _04363_
+ sg13g2_a22oi_1
X_24086_ _03987_ VPWR VGND _04364_ sg13g2_buf_1
X_24087_ _03827_ VPWR VGND _04365_ sg13g2_buf_1
X_24088_ _02147_ _03822_ VPWR VGND _04366_ sg13g2_nand2b_1
X_24089_ _04365_ _02171_ _04366_ VPWR VGND _04367_ sg13g2_o21ai_1
X_24090_ _04364_ _04367_ _03740_ VPWR VGND _04368_ sg13g2_a21oi_1
X_24091_ _04355_ _04363_ _04368_ VPWR VGND _04369_ sg13g2_a21oi_1
X_24092_ _00145_ _04353_ _04354_ _02210_ _04369_ VPWR 
+ VGND
+ _04370_ sg13g2_a221oi_1
X_24093_ _03720_ VPWR VGND _04371_ sg13g2_buf_1
X_24094_ _04075_ VPWR VGND _04372_ sg13g2_buf_1
X_24095_ _04372_ VPWR VGND _04373_ sg13g2_buf_1
X_24096_ _00143_ _03969_ VPWR VGND _04374_ sg13g2_nand2_1
X_24097_ \atbs_core_0.spike_memory_0.n2409_o[11]\ _04373_ _04374_ VPWR VGND _04375_ sg13g2_o21ai_1
X_24098_ _04002_ VPWR VGND _04376_ sg13g2_buf_1
X_24099_ _04376_ VPWR VGND _04377_ sg13g2_buf_1
X_24100_ _03744_ VPWR VGND _04378_ sg13g2_buf_1
X_24101_ _03761_ VPWR VGND _04379_ sg13g2_buf_1
X_24102_ _04379_ _02630_ VPWR VGND _04380_ sg13g2_nor2_1
X_24103_ _04280_ VPWR VGND _04381_ sg13g2_buf_1
X_24104_ _02651_ _04381_ VPWR VGND _04382_ sg13g2_nor2_1
X_24105_ _03978_ VPWR VGND _04383_ sg13g2_buf_1
X_24106_ _04383_ VPWR VGND _04384_ sg13g2_buf_1
X_24107_ _04378_ _04380_ _04382_ _04384_ VPWR VGND 
+ _04385_
+ sg13g2_a22oi_1
X_24108_ _04009_ VPWR VGND _04386_ sg13g2_buf_1
X_24109_ _04386_ VPWR VGND _04387_ sg13g2_buf_1
X_24110_ _04387_ VPWR VGND _04388_ sg13g2_buf_1
X_24111_ _02630_ _04268_ VPWR VGND _04389_ sg13g2_nand2b_1
X_24112_ _04383_ _02651_ _04389_ VPWR VGND _04390_ sg13g2_o21ai_1
X_24113_ _03767_ VPWR VGND _04391_ sg13g2_buf_1
X_24114_ _04391_ VPWR VGND _04392_ sg13g2_buf_1
X_24115_ _04392_ VPWR VGND _04393_ sg13g2_buf_1
X_24116_ _04388_ _04390_ _04393_ VPWR VGND _04394_ sg13g2_a21oi_1
X_24117_ _04377_ _04385_ _04394_ VPWR VGND _04395_ sg13g2_a21oi_1
X_24118_ _12079_ _04375_ _04395_ VPWR VGND _04396_ sg13g2_nor3_1
X_24119_ _04337_ _04352_ _04370_ _04371_ _04396_ VPWR 
+ VGND
+ _04397_ sg13g2_a221oi_1
X_24120_ \atbs_core_0.spike_memory_0.n2413_o[11]\ _03776_ VPWR VGND _04398_ sg13g2_nor2_1
X_24121_ \atbs_core_0.spike_memory_0.n2410_o[11]\ _03806_ VPWR VGND _04399_ sg13g2_nor2_1
X_24122_ _03855_ _12530_ VPWR VGND _04400_ sg13g2_nor2_1
X_24123_ _12553_ _03951_ VPWR VGND _04401_ sg13g2_nor2_1
X_24124_ _04047_ _04400_ _04401_ _04052_ VPWR VGND 
+ _04402_
+ sg13g2_a22oi_1
X_24125_ _12530_ _04054_ VPWR VGND _04403_ sg13g2_nand2b_1
X_24126_ _04051_ _12553_ _04403_ VPWR VGND _04404_ sg13g2_o21ai_1
X_24127_ _03955_ _04404_ _03868_ VPWR VGND _04405_ sg13g2_a21oi_1
X_24128_ _03993_ _04402_ _04405_ VPWR VGND _04406_ sg13g2_a21oi_1
X_24129_ _03800_ _04398_ _04399_ _04406_ VPWR VGND 
+ _04407_
+ sg13g2_nor4_1
X_24130_ \atbs_core_0.spike_memory_0.n2417_o[11]\ _04076_ VPWR VGND _04408_ sg13g2_nor2_1
X_24131_ \atbs_core_0.spike_memory_0.n2414_o[11]\ _03806_ _03723_ VPWR VGND _04409_ sg13g2_o21ai_1
X_24132_ _04089_ _12585_ VPWR VGND _04410_ sg13g2_nor2_1
X_24133_ _12608_ _04086_ VPWR VGND _04411_ sg13g2_nor2_1
X_24134_ _04082_ _04410_ _04411_ _04090_ VPWR VGND 
+ _04412_
+ sg13g2_a22oi_1
X_24135_ _04011_ VPWR VGND _04413_ sg13g2_buf_1
X_24136_ _12585_ _04094_ VPWR VGND _04414_ sg13g2_nand2b_1
X_24137_ _04413_ _12608_ _04414_ VPWR VGND _04415_ sg13g2_o21ai_1
X_24138_ _04092_ _04415_ _04098_ VPWR VGND _04416_ sg13g2_a21oi_1
X_24139_ _04081_ _04412_ _04416_ VPWR VGND _04417_ sg13g2_a21oi_1
X_24140_ _04408_ _04409_ _04417_ VPWR VGND _04418_ sg13g2_nor3_1
X_24141_ \atbs_core_0.spike_memory_0.n2436_q[1208]\ _04245_ VPWR VGND _04419_ sg13g2_nor2_1
X_24142_ \atbs_core_0.spike_memory_0.n2418_o[11]\ _04247_ VPWR VGND _04420_ sg13g2_nor2_1
X_24143_ _03989_ _12644_ VPWR VGND _04421_ sg13g2_nor2_1
X_24144_ _04085_ VPWR VGND _04422_ sg13g2_buf_1
X_24145_ _12667_ _04422_ VPWR VGND _04423_ sg13g2_nor2_1
X_24146_ _04280_ _04421_ _04423_ _04283_ VPWR VGND 
+ _04424_
+ sg13g2_a22oi_1
X_24147_ _04093_ VPWR VGND _04425_ sg13g2_buf_1
X_24148_ _12644_ _04425_ VPWR VGND _04426_ sg13g2_nand2b_1
X_24149_ _03847_ _12667_ _04426_ VPWR VGND _04427_ sg13g2_o21ai_1
X_24150_ _03860_ _04427_ _04287_ VPWR VGND _04428_ sg13g2_a21oi_1
X_24151_ _04392_ _04424_ _04428_ VPWR VGND _04429_ sg13g2_a21oi_1
X_24152_ _12094_ _04419_ _04420_ _04429_ VPWR VGND 
+ _04430_
+ sg13g2_nor4_1
X_24153_ _04407_ _04418_ _04430_ VPWR VGND _04431_ sg13g2_nor3_1
X_24154_ \atbs_core_0.spike_memory_0.n2385_o[11]\ _03970_ VPWR VGND _04432_ sg13g2_nand2b_1
X_24155_ \atbs_core_0.spike_memory_0.n2382_o[11]\ _04292_ _04432_ VPWR VGND _04433_ sg13g2_o21ai_1
X_24156_ _04011_ _02299_ VPWR VGND _04434_ sg13g2_nor2_1
X_24157_ _02324_ _04107_ VPWR VGND _04435_ sg13g2_nor2_1
X_24158_ _03750_ _04434_ _04435_ _04413_ VPWR VGND 
+ _04436_
+ sg13g2_a22oi_1
X_24159_ _02299_ _04093_ VPWR VGND _04437_ sg13g2_nand2b_1
X_24160_ _04088_ _02324_ _04437_ VPWR VGND _04438_ sg13g2_o21ai_1
X_24161_ _03986_ _04438_ _04097_ VPWR VGND _04439_ sg13g2_a21oi_1
X_24162_ _03768_ _04436_ _04439_ VPWR VGND _04440_ sg13g2_a21oi_1
X_24163_ _04433_ _04440_ VPWR VGND _04441_ sg13g2_or2_1
X_24164_ _12084_ VPWR VGND _04442_ sg13g2_buf_1
X_24165_ \atbs_core_0.spike_memory_0.n2381_o[11]\ _04442_ VPWR VGND _04443_ sg13g2_nor2_1
X_24166_ \atbs_core_0.spike_memory_0.n2378_o[11]\ _03999_ VPWR VGND _04444_ sg13g2_nor2_1
X_24167_ _03890_ _02245_ VPWR VGND _04445_ sg13g2_nor2_1
X_24168_ _02267_ _03741_ VPWR VGND _04446_ sg13g2_nor2_1
X_24169_ _03850_ _04445_ _04446_ _03791_ VPWR VGND 
+ _04447_
+ sg13g2_a22oi_1
X_24170_ _02245_ _03845_ VPWR VGND _04448_ sg13g2_nand2b_1
X_24171_ _03890_ _02267_ _04448_ VPWR VGND _04449_ sg13g2_o21ai_1
X_24172_ _03730_ _04449_ _03809_ VPWR VGND _04450_ sg13g2_a21oi_1
X_24173_ _03867_ _04447_ _04450_ VPWR VGND _04451_ sg13g2_a21oi_1
X_24174_ _03726_ _04443_ _04444_ _04451_ VPWR VGND 
+ _04452_
+ sg13g2_nor4_1
X_24175_ \atbs_core_0.spike_memory_0.n2389_o[11]\ _04442_ VPWR VGND _04453_ sg13g2_nor2_1
X_24176_ \atbs_core_0.spike_memory_0.n2386_o[11]\ _03999_ VPWR VGND _04454_ sg13g2_nor2_1
X_24177_ _02709_ VPWR VGND _04455_ sg13g2_buf_1
X_24178_ _04455_ _02355_ VPWR VGND _04456_ sg13g2_nor2_1
X_24179_ _02378_ _03741_ VPWR VGND _04457_ sg13g2_nor2_1
X_24180_ _04085_ _04456_ _04457_ _03915_ VPWR VGND 
+ _04458_
+ sg13g2_a22oi_1
X_24181_ _02355_ _03845_ VPWR VGND _04459_ sg13g2_nand2b_1
X_24182_ _04455_ _02378_ _04459_ VPWR VGND _04460_ sg13g2_o21ai_1
X_24183_ _04009_ _04460_ _03809_ VPWR VGND _04461_ sg13g2_a21oi_1
X_24184_ _04068_ _04458_ _04461_ VPWR VGND _04462_ sg13g2_a21oi_1
X_24185_ _07555_ _04453_ _04454_ _04462_ VPWR VGND 
+ _04463_
+ sg13g2_nor4_1
X_24186_ _04452_ _04463_ _12090_ VPWR VGND _04464_ sg13g2_o21ai_1
X_24187_ _04276_ _04441_ _04464_ VPWR VGND _04465_ sg13g2_o21ai_1
X_24188_ \atbs_core_0.spike_memory_0.n2401_o[11]\ _03970_ VPWR VGND _04466_ sg13g2_nand2b_1
X_24189_ \atbs_core_0.spike_memory_0.n2398_o[11]\ _04078_ _04466_ VPWR VGND _04467_ sg13g2_o21ai_1
X_24190_ _03891_ _02535_ VPWR VGND _04468_ sg13g2_nor2_1
X_24191_ _02556_ _04107_ VPWR VGND _04469_ sg13g2_nor2_1
X_24192_ _03818_ _04468_ _04469_ _04346_ VPWR VGND 
+ _04470_
+ sg13g2_a22oi_1
X_24193_ _02535_ _02710_ VPWR VGND _04471_ sg13g2_nand2b_1
X_24194_ _03763_ _02556_ _04471_ VPWR VGND _04472_ sg13g2_o21ai_1
X_24195_ _03986_ _04472_ _02699_ VPWR VGND _04473_ sg13g2_a21oi_1
X_24196_ _03830_ _04470_ _04473_ VPWR VGND _04474_ sg13g2_a21oi_1
X_24197_ _04467_ _04474_ VPWR VGND _04475_ sg13g2_or2_1
X_24198_ \atbs_core_0.spike_memory_0.n2397_o[11]\ _04442_ VPWR VGND _04476_ sg13g2_nor2_1
X_24199_ \atbs_core_0.spike_memory_0.n2394_o[11]\ _03999_ VPWR VGND _04477_ sg13g2_nor2_1
X_24200_ _03862_ _02488_ VPWR VGND _04478_ sg13g2_nor2_1
X_24201_ _02509_ _03749_ VPWR VGND _04479_ sg13g2_nor2_1
X_24202_ _03862_ VPWR VGND _04480_ sg13g2_buf_1
X_24203_ _04085_ _04478_ _04479_ _04480_ VPWR VGND 
+ _04481_
+ sg13g2_a22oi_1
X_24204_ _02488_ _03845_ VPWR VGND _04482_ sg13g2_nand2b_1
X_24205_ _03862_ _02509_ _04482_ VPWR VGND _04483_ sg13g2_o21ai_1
X_24206_ _04009_ _04483_ _03809_ VPWR VGND _04484_ sg13g2_a21oi_1
X_24207_ _04097_ _04481_ _04484_ VPWR VGND _04485_ sg13g2_a21oi_1
X_24208_ _03726_ _04476_ _04477_ _04485_ VPWR VGND 
+ _04486_
+ sg13g2_nor4_1
X_24209_ \atbs_core_0.spike_memory_0.n2405_o[11]\ _04442_ VPWR VGND _04487_ sg13g2_nor2_1
X_24210_ \atbs_core_0.spike_memory_0.n2402_o[11]\ _03778_ VPWR VGND _04488_ sg13g2_nor2_1
X_24211_ _04093_ _02583_ VPWR VGND _04489_ sg13g2_nor2_1
X_24212_ _02604_ _03749_ VPWR VGND _04490_ sg13g2_nor2_1
X_24213_ _04107_ _04489_ _04490_ _03982_ VPWR VGND 
+ _04491_
+ sg13g2_a22oi_1
X_24214_ _02583_ _03762_ VPWR VGND _04492_ sg13g2_nand2b_1
X_24215_ _03981_ _02604_ _04492_ VPWR VGND _04493_ sg13g2_o21ai_1
X_24216_ _04009_ _04493_ _03809_ VPWR VGND _04494_ sg13g2_a21oi_1
X_24217_ _02699_ _04491_ _04494_ VPWR VGND _04495_ sg13g2_a21oi_1
X_24218_ _07555_ _04487_ _04488_ _04495_ VPWR VGND 
+ _04496_
+ sg13g2_nor4_1
X_24219_ _04486_ _04496_ _12090_ VPWR VGND _04497_ sg13g2_o21ai_1
X_24220_ _03924_ _04475_ _04497_ VPWR VGND _04498_ sg13g2_o21ai_1
X_24221_ _07547_ _04465_ _04498_ _03717_ VPWR VGND 
+ _04499_
+ sg13g2_a22oi_1
X_24222_ _12079_ _04431_ _04499_ VPWR VGND _04500_ sg13g2_o21ai_1
X_24223_ _04336_ _04500_ VPWR VGND _04501_ sg13g2_nor2_1
X_24224_ _04336_ _04397_ _04501_ VPWR VGND _04502_ sg13g2_a21oi_1
X_24225_ _07549_ VPWR VGND _04503_ sg13g2_buf_1
X_24226_ _03925_ VPWR VGND _04504_ sg13g2_buf_1
X_24227_ _03774_ VPWR VGND _04505_ sg13g2_buf_1
X_24228_ _04372_ VPWR VGND _04506_ sg13g2_buf_1
X_24229_ \atbs_core_0.spike_memory_0.n2361_o[11]\ _04506_ VPWR VGND _04507_ sg13g2_nor2_1
X_24230_ _04032_ VPWR VGND _04508_ sg13g2_buf_1
X_24231_ \atbs_core_0.spike_memory_0.n2358_o[11]\ _04508_ VPWR VGND _04509_ sg13g2_nor2_1
X_24232_ _04003_ VPWR VGND _04510_ sg13g2_buf_1
X_24233_ _04510_ VPWR VGND _04511_ sg13g2_buf_1
X_24234_ _04237_ VPWR VGND _04512_ sg13g2_buf_1
X_24235_ _04512_ VPWR VGND _04513_ sg13g2_buf_1
X_24236_ _04513_ _02131_ VPWR VGND _04514_ sg13g2_nor2_1
X_24237_ _02316_ _04381_ VPWR VGND _04515_ sg13g2_nor2_1
X_24238_ _04511_ _04514_ _04515_ _04384_ VPWR VGND 
+ _04516_
+ sg13g2_a22oi_1
X_24239_ _04387_ VPWR VGND _04517_ sg13g2_buf_1
X_24240_ _04267_ VPWR VGND _04518_ sg13g2_buf_1
X_24241_ _02131_ _04518_ VPWR VGND _04519_ sg13g2_nand2b_1
X_24242_ _04383_ _02316_ _04519_ VPWR VGND _04520_ sg13g2_o21ai_1
X_24243_ _03840_ VPWR VGND _04521_ sg13g2_buf_1
X_24244_ _04517_ _04520_ _04521_ VPWR VGND _04522_ sg13g2_a21oi_1
X_24245_ _04377_ _04516_ _04522_ VPWR VGND _04523_ sg13g2_a21oi_1
X_24246_ _04505_ _04507_ _04509_ _04523_ VPWR VGND 
+ _04524_
+ sg13g2_nor4_1
X_24247_ _03877_ VPWR VGND _04525_ sg13g2_buf_1
X_24248_ \atbs_core_0.spike_memory_0.n2369_o[11]\ _04525_ VPWR VGND _04526_ sg13g2_nor2_1
X_24249_ _03835_ VPWR VGND _04527_ sg13g2_buf_1
X_24250_ _04527_ VPWR VGND _04528_ sg13g2_buf_1
X_24251_ \atbs_core_0.spike_memory_0.n2366_o[11]\ _04528_ VPWR VGND _04529_ sg13g2_nor2_1
X_24252_ _04021_ VPWR VGND _04530_ sg13g2_buf_1
X_24253_ _04359_ VPWR VGND _04531_ sg13g2_buf_1
X_24254_ _03887_ _02038_ VPWR VGND _04532_ sg13g2_nor2_1
X_24255_ _04023_ VPWR VGND _04533_ sg13g2_buf_1
X_24256_ _02060_ _04533_ VPWR VGND _04534_ sg13g2_nor2_1
X_24257_ _03761_ VPWR VGND _04535_ sg13g2_buf_1
X_24258_ _04535_ VPWR VGND _04536_ sg13g2_buf_1
X_24259_ _04531_ _04532_ _04534_ _04536_ VPWR VGND 
+ _04537_
+ sg13g2_a22oi_1
X_24260_ _03759_ VPWR VGND _04538_ sg13g2_buf_1
X_24261_ _03747_ VPWR VGND _04539_ sg13g2_buf_1
X_24262_ _02038_ _04347_ VPWR VGND _04540_ sg13g2_nand2b_1
X_24263_ _04539_ _02060_ _04540_ VPWR VGND _04541_ sg13g2_o21ai_1
X_24264_ _04081_ VPWR VGND _04542_ sg13g2_buf_1
X_24265_ _04538_ _04541_ _04542_ VPWR VGND _04543_ sg13g2_a21oi_1
X_24266_ _04530_ _04537_ _04543_ VPWR VGND _04544_ sg13g2_a21oi_1
X_24267_ _04126_ _04526_ _04529_ _04544_ VPWR VGND 
+ _04545_
+ sg13g2_nor4_1
X_24268_ _04504_ _04524_ _04545_ VPWR VGND _04546_ sg13g2_nor3_1
X_24269_ _03724_ VPWR VGND _04547_ sg13g2_buf_1
X_24270_ \atbs_core_0.spike_memory_0.n2365_o[11]\ _04525_ VPWR VGND _04548_ sg13g2_nor2_1
X_24271_ _04527_ VPWR VGND _04549_ sg13g2_buf_1
X_24272_ \atbs_core_0.spike_memory_0.n2362_o[11]\ _04549_ VPWR VGND _04550_ sg13g2_nor2_1
X_24273_ _04021_ VPWR VGND _04551_ sg13g2_buf_1
X_24274_ _02711_ VPWR VGND _04552_ sg13g2_buf_1
X_24275_ _04552_ VPWR VGND _04553_ sg13g2_buf_1
X_24276_ _04553_ _12568_ VPWR VGND _04554_ sg13g2_nor2_1
X_24277_ _04082_ VPWR VGND _04555_ sg13g2_buf_1
X_24278_ _02011_ _04555_ VPWR VGND _04556_ sg13g2_nor2_1
X_24279_ _04535_ VPWR VGND _04557_ sg13g2_buf_1
X_24280_ _04378_ _04554_ _04556_ _04557_ VPWR VGND 
+ _04558_
+ sg13g2_a22oi_1
X_24281_ _04105_ VPWR VGND _04559_ sg13g2_buf_1
X_24282_ _12568_ _04559_ VPWR VGND _04560_ sg13g2_nand2b_1
X_24283_ _03755_ _02011_ _04560_ VPWR VGND _04561_ sg13g2_o21ai_1
X_24284_ _04081_ VPWR VGND _04562_ sg13g2_buf_1
X_24285_ _04388_ _04561_ _04562_ VPWR VGND _04563_ sg13g2_a21oi_1
X_24286_ _04551_ _04558_ _04563_ VPWR VGND _04564_ sg13g2_a21oi_1
X_24287_ _03729_ _04548_ _04550_ _04564_ VPWR VGND 
+ _04565_
+ sg13g2_nor4_1
X_24288_ \atbs_core_0.spike_memory_0.n2373_o[11]\ _12088_ VPWR VGND _04566_ sg13g2_nor2_1
X_24289_ \atbs_core_0.spike_memory_0.n2370_o[11]\ _04528_ VPWR VGND _04567_ sg13g2_nor2_1
X_24290_ _03929_ VPWR VGND _04568_ sg13g2_buf_1
X_24291_ _03934_ _02092_ VPWR VGND _04569_ sg13g2_nor2_1
X_24292_ _03884_ VPWR VGND _04570_ sg13g2_buf_1
X_24293_ _02115_ _04570_ VPWR VGND _04571_ sg13g2_nor2_1
X_24294_ _04568_ _04569_ _04571_ _02714_ VPWR VGND 
+ _04572_
+ sg13g2_a22oi_1
X_24295_ _03889_ VPWR VGND _04573_ sg13g2_buf_1
X_24296_ _03882_ VPWR VGND _04574_ sg13g2_buf_1
X_24297_ _02092_ _04361_ VPWR VGND _04575_ sg13g2_nand2b_1
X_24298_ _04574_ _02115_ _04575_ VPWR VGND _04576_ sg13g2_o21ai_1
X_24299_ _04573_ _04576_ _04338_ VPWR VGND _04577_ sg13g2_a21oi_1
X_24300_ _02702_ _04572_ _04577_ VPWR VGND _04578_ sg13g2_a21oi_1
X_24301_ _04126_ _04566_ _04567_ _04578_ VPWR VGND 
+ _04579_
+ sg13g2_nor4_1
X_24302_ _04547_ _04565_ _04579_ VPWR VGND _04580_ sg13g2_nor3_1
X_24303_ _04503_ _04546_ _04580_ VPWR VGND _04581_ sg13g2_nor3_1
X_24304_ _04333_ _04502_ _04581_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[11]\ sg13g2_a21o_1
X_24305_ _04372_ VPWR VGND _04582_ sg13g2_buf_1
X_24306_ \atbs_core_0.spike_memory_0.n2365_o[12]\ _04582_ VPWR VGND _04583_ sg13g2_nor2_1
X_24307_ _04230_ VPWR VGND _04584_ sg13g2_buf_1
X_24308_ \atbs_core_0.spike_memory_0.n2362_o[12]\ _04584_ VPWR VGND _04585_ sg13g2_nor2_1
X_24309_ _03869_ VPWR VGND _04586_ sg13g2_buf_1
X_24310_ _03851_ VPWR VGND _04587_ sg13g2_buf_1
X_24311_ _04587_ VPWR VGND _04588_ sg13g2_buf_1
X_24312_ _03863_ VPWR VGND _04589_ sg13g2_buf_1
X_24313_ _04589_ VPWR VGND _04590_ sg13g2_buf_1
X_24314_ _04590_ _12571_ VPWR VGND _04591_ sg13g2_nor2_1
X_24315_ _02012_ _04150_ VPWR VGND _04592_ sg13g2_nor2_1
X_24316_ _04167_ VPWR VGND _04593_ sg13g2_buf_1
X_24317_ _04593_ VPWR VGND _04594_ sg13g2_buf_1
X_24318_ _04588_ _04591_ _04592_ _04594_ VPWR VGND 
+ _04595_
+ sg13g2_a22oi_1
X_24319_ _03987_ VPWR VGND _04596_ sg13g2_buf_1
X_24320_ _03846_ VPWR VGND _04597_ sg13g2_buf_1
X_24321_ _04597_ VPWR VGND _04598_ sg13g2_buf_1
X_24322_ _12571_ _04598_ VPWR VGND _04599_ sg13g2_nand2b_1
X_24323_ _04593_ _02012_ _04599_ VPWR VGND _04600_ sg13g2_o21ai_1
X_24324_ _04596_ _04600_ _02701_ VPWR VGND _04601_ sg13g2_a21oi_1
X_24325_ _04586_ _04595_ _04601_ VPWR VGND _04602_ sg13g2_a21oi_1
X_24326_ _04505_ _04583_ _04585_ _04602_ VPWR VGND 
+ _04603_
+ sg13g2_nor4_1
X_24327_ _03900_ VPWR VGND _04604_ sg13g2_buf_1
X_24328_ \atbs_core_0.spike_memory_0.n2373_o[12]\ _04373_ VPWR VGND _04605_ sg13g2_nor2_1
X_24329_ _04230_ VPWR VGND _04606_ sg13g2_buf_1
X_24330_ \atbs_core_0.spike_memory_0.n2370_o[12]\ _04606_ VPWR VGND _04607_ sg13g2_nor2_1
X_24331_ _03974_ VPWR VGND _04608_ sg13g2_buf_1
X_24332_ _04587_ VPWR VGND _04609_ sg13g2_buf_1
X_24333_ _04589_ VPWR VGND _04610_ sg13g2_buf_1
X_24334_ _04610_ _02093_ VPWR VGND _04611_ sg13g2_nor2_1
X_24335_ _02116_ _03814_ VPWR VGND _04612_ sg13g2_nor2_1
X_24336_ _04610_ VPWR VGND _04613_ sg13g2_buf_1
X_24337_ _04609_ _04611_ _04612_ _04613_ VPWR VGND 
+ _04614_
+ sg13g2_a22oi_1
X_24338_ _03987_ VPWR VGND _04615_ sg13g2_buf_1
X_24339_ _04589_ VPWR VGND _04616_ sg13g2_buf_1
X_24340_ _02093_ _04283_ VPWR VGND _04617_ sg13g2_nand2b_1
X_24341_ _04616_ _02116_ _04617_ VPWR VGND _04618_ sg13g2_o21ai_1
X_24342_ _04615_ _04618_ _03948_ VPWR VGND _04619_ sg13g2_a21oi_1
X_24343_ _04608_ _04614_ _04619_ VPWR VGND _04620_ sg13g2_a21oi_1
X_24344_ _04604_ _04605_ _04607_ _04620_ VPWR VGND 
+ _04621_
+ sg13g2_nor4_1
X_24345_ _04603_ _04621_ _04504_ VPWR VGND _04622_ sg13g2_o21ai_1
X_24346_ _04245_ VPWR VGND _04623_ sg13g2_buf_1
X_24347_ \atbs_core_0.spike_memory_0.n2361_o[12]\ _04623_ VPWR VGND _04624_ sg13g2_nor2_1
X_24348_ \atbs_core_0.spike_memory_0.n2358_o[12]\ _04584_ VPWR VGND _04625_ sg13g2_nor2_1
X_24349_ _03869_ VPWR VGND _04626_ sg13g2_buf_1
X_24350_ _04593_ _02133_ VPWR VGND _04627_ sg13g2_nor2_1
X_24351_ _03782_ VPWR VGND _04628_ sg13g2_buf_1
X_24352_ _02329_ _04628_ VPWR VGND _04629_ sg13g2_nor2_1
X_24353_ _04357_ VPWR VGND _04630_ sg13g2_buf_1
X_24354_ _04588_ _04627_ _04629_ _04630_ VPWR VGND 
+ _04631_
+ sg13g2_a22oi_1
X_24355_ _04167_ VPWR VGND _04632_ sg13g2_buf_1
X_24356_ _02133_ _04052_ VPWR VGND _04633_ sg13g2_nand2b_1
X_24357_ _04632_ _02329_ _04633_ VPWR VGND _04634_ sg13g2_o21ai_1
X_24358_ _02700_ VPWR VGND _04635_ sg13g2_buf_1
X_24359_ _04596_ _04634_ _04635_ VPWR VGND _04636_ sg13g2_a21oi_1
X_24360_ _04626_ _04631_ _04636_ VPWR VGND _04637_ sg13g2_a21oi_1
X_24361_ _03872_ _04624_ _04625_ _04637_ VPWR VGND 
+ _04638_
+ sg13g2_nor4_1
X_24362_ \atbs_core_0.spike_memory_0.n2369_o[12]\ _04582_ VPWR VGND _04639_ sg13g2_nor2_1
X_24363_ \atbs_core_0.spike_memory_0.n2366_o[12]\ _04606_ VPWR VGND _04640_ sg13g2_nor2_1
X_24364_ _04616_ _02039_ VPWR VGND _04641_ sg13g2_nor2_1
X_24365_ _02061_ _04035_ VPWR VGND _04642_ sg13g2_nor2_1
X_24366_ _04609_ _04641_ _04642_ _04594_ VPWR VGND 
+ _04643_
+ sg13g2_a22oi_1
X_24367_ _02039_ _03848_ VPWR VGND _04644_ sg13g2_nand2b_1
X_24368_ _04590_ _02061_ _04644_ VPWR VGND _04645_ sg13g2_o21ai_1
X_24369_ _04615_ _04645_ _04149_ VPWR VGND _04646_ sg13g2_a21oi_1
X_24370_ _04586_ _04643_ _04646_ VPWR VGND _04647_ sg13g2_a21oi_1
X_24371_ _04219_ _04639_ _04640_ _04647_ VPWR VGND 
+ _04648_
+ sg13g2_nor4_1
X_24372_ _04638_ _04648_ _04547_ VPWR VGND _04649_ sg13g2_o21ai_1
X_24373_ _04622_ _04649_ VPWR VGND _04650_ sg13g2_and2_1
X_24374_ _03937_ VPWR VGND _04651_ sg13g2_buf_1
X_24375_ _04651_ _02403_ VPWR VGND _04652_ sg13g2_nor2_1
X_24376_ _02422_ _04510_ VPWR VGND _04653_ sg13g2_nor2_1
X_24377_ _04356_ _04652_ _04653_ _04362_ VPWR VGND 
+ _04654_
+ sg13g2_a22oi_1
X_24378_ _02403_ _03882_ VPWR VGND _04655_ sg13g2_nand2b_1
X_24379_ _04320_ _02422_ _04655_ VPWR VGND _04656_ sg13g2_o21ai_1
X_24380_ _04364_ _04656_ _04376_ VPWR VGND _04657_ sg13g2_a21oi_1
X_24381_ _04355_ _04654_ _04657_ VPWR VGND _04658_ sg13g2_a21oi_1
X_24382_ _00147_ _04353_ _04354_ _02457_ _04658_ VPWR 
+ VGND
+ _04659_ sg13g2_a221oi_1
X_24383_ _03732_ VPWR VGND _04660_ sg13g2_buf_1
X_24384_ _03972_ VPWR VGND _04661_ sg13g2_buf_1
X_24385_ _04587_ VPWR VGND _04662_ sg13g2_buf_1
X_24386_ _04632_ _02631_ VPWR VGND _04663_ sg13g2_nor2_1
X_24387_ _02652_ _04628_ VPWR VGND _04664_ sg13g2_nor2_1
X_24388_ _04662_ _04663_ _04664_ _04630_ VPWR VGND 
+ _04665_
+ sg13g2_a22oi_1
X_24389_ _03987_ VPWR VGND _04666_ sg13g2_buf_1
X_24390_ _02631_ _03957_ VPWR VGND _04667_ sg13g2_nand2b_1
X_24391_ _04357_ _02652_ _04667_ VPWR VGND _04668_ sg13g2_o21ai_1
X_24392_ _04666_ _04668_ _03880_ VPWR VGND _04669_ sg13g2_a21oi_1
X_24393_ _04626_ _04665_ _04669_ VPWR VGND _04670_ sg13g2_a21oi_1
X_24394_ _00146_ _04660_ _04661_ _02682_ _04670_ VPWR 
+ VGND
+ _04671_ sg13g2_a221oi_1
X_24395_ _07541_ _07547_ VPWR VGND _04672_ sg13g2_nor2_1
X_24396_ _04672_ VPWR VGND _04673_ sg13g2_buf_1
X_24397_ _03718_ _04659_ _04671_ _04673_ VPWR VGND 
+ _04674_
+ sg13g2_a22oi_1
X_24398_ _03732_ VPWR VGND _04675_ sg13g2_buf_1
X_24399_ _03736_ VPWR VGND _04676_ sg13g2_buf_1
X_24400_ _03831_ VPWR VGND _04677_ sg13g2_buf_1
X_24401_ _04651_ _02149_ VPWR VGND _04678_ sg13g2_nor2_1
X_24402_ _02172_ _04510_ VPWR VGND _04679_ sg13g2_nor2_1
X_24403_ _04347_ VPWR VGND _04680_ sg13g2_buf_1
X_24404_ _04339_ _04678_ _04679_ _04680_ VPWR VGND 
+ _04681_
+ sg13g2_a22oi_1
X_24405_ _02149_ _04552_ VPWR VGND _04682_ sg13g2_nand2b_1
X_24406_ _04340_ _02172_ _04682_ VPWR VGND _04683_ sg13g2_o21ai_1
X_24407_ _04002_ VPWR VGND _04684_ sg13g2_buf_1
X_24408_ _04345_ _04683_ _04684_ VPWR VGND _04685_ sg13g2_a21oi_1
X_24409_ _04677_ _04681_ _04685_ VPWR VGND _04686_ sg13g2_a21oi_1
X_24410_ _00148_ _04675_ _04676_ _02212_ _04686_ VPWR 
+ VGND
+ _04687_ sg13g2_a221oi_1
X_24411_ _07556_ VPWR VGND _04688_ sg13g2_buf_1
X_24412_ _04371_ _04687_ _04688_ VPWR VGND _04689_ sg13g2_a21oi_1
X_24413_ _04674_ _04689_ VPWR VGND _04690_ sg13g2_nand2_1
X_24414_ \atbs_core_0.spike_memory_0.n2413_o[12]\ _03901_ VPWR VGND _04691_ sg13g2_nor2_1
X_24415_ \atbs_core_0.spike_memory_0.n2410_o[12]\ _03807_ VPWR VGND _04692_ sg13g2_nor2_1
X_24416_ _03816_ _12531_ VPWR VGND _04693_ sg13g2_nor2_1
X_24417_ _12554_ _03819_ VPWR VGND _04694_ sg13g2_nor2_1
X_24418_ _04035_ _04693_ _04694_ _03823_ VPWR VGND 
+ _04695_
+ sg13g2_a22oi_1
X_24419_ _12531_ _03916_ VPWR VGND _04696_ sg13g2_nand2b_1
X_24420_ _03930_ _12554_ _04696_ VPWR VGND _04697_ sg13g2_o21ai_1
X_24421_ _03825_ _04697_ _03831_ VPWR VGND _04698_ sg13g2_a21oi_1
X_24422_ _03812_ _04695_ _04698_ VPWR VGND _04699_ sg13g2_a21oi_1
X_24423_ _04074_ _04691_ _04692_ _04699_ VPWR VGND 
+ _04700_
+ sg13g2_nor4_1
X_24424_ \atbs_core_0.spike_memory_0.n2417_o[12]\ _04623_ VPWR VGND _04701_ sg13g2_nor2_1
X_24425_ _03835_ VPWR VGND _04702_ sg13g2_buf_1
X_24426_ \atbs_core_0.spike_memory_0.n2414_o[12]\ _04702_ _03966_ VPWR VGND _04703_ sg13g2_o21ai_1
X_24427_ _03989_ VPWR VGND _04704_ sg13g2_buf_1
X_24428_ _04704_ _12586_ VPWR VGND _04705_ sg13g2_nor2_1
X_24429_ _12610_ _04587_ VPWR VGND _04706_ sg13g2_nor2_1
X_24430_ _04381_ _04705_ _04706_ _04343_ VPWR VGND 
+ _04707_
+ sg13g2_a22oi_1
X_24431_ _03847_ VPWR VGND _04708_ sg13g2_buf_1
X_24432_ _12586_ _04589_ VPWR VGND _04709_ sg13g2_nand2b_1
X_24433_ _04708_ _12610_ _04709_ VPWR VGND _04710_ sg13g2_o21ai_1
X_24434_ _03861_ _04710_ _03869_ VPWR VGND _04711_ sg13g2_a21oi_1
X_24435_ _04393_ _04707_ _04711_ VPWR VGND _04712_ sg13g2_a21oi_1
X_24436_ _04701_ _04703_ _04712_ VPWR VGND _04713_ sg13g2_nor3_1
X_24437_ \atbs_core_0.spike_memory_0.n2436_q[1209]\ _03804_ VPWR VGND _04714_ sg13g2_nor2_1
X_24438_ \atbs_core_0.spike_memory_0.n2418_o[12]\ _03946_ VPWR VGND _04715_ sg13g2_nor2_1
X_24439_ _03843_ VPWR VGND _04716_ sg13g2_buf_1
X_24440_ _03848_ _12645_ VPWR VGND _04717_ sg13g2_nor2_1
X_24441_ _12670_ _03852_ VPWR VGND _04718_ sg13g2_nor2_1
X_24442_ _04716_ _04717_ _04718_ _03857_ VPWR VGND 
+ _04719_
+ sg13g2_a22oi_1
X_24443_ _12645_ _03864_ VPWR VGND _04720_ sg13g2_nand2b_1
X_24444_ _04598_ _12670_ _04720_ VPWR VGND _04721_ sg13g2_o21ai_1
X_24445_ _03861_ _04721_ _03869_ VPWR VGND _04722_ sg13g2_a21oi_1
X_24446_ _03841_ _04719_ _04722_ VPWR VGND _04723_ sg13g2_a21oi_1
X_24447_ _12095_ _04714_ _04715_ _04723_ VPWR VGND 
+ _04724_
+ sg13g2_nor4_1
X_24448_ _04700_ _04713_ _04724_ VPWR VGND _04725_ sg13g2_nor3_1
X_24449_ \atbs_core_0.spike_memory_0.n2385_o[12]\ _03735_ VPWR VGND _04726_ sg13g2_nand2b_1
X_24450_ \atbs_core_0.spike_memory_0.n2382_o[12]\ _03779_ _04726_ VPWR VGND _04727_ sg13g2_o21ai_1
X_24451_ _03746_ _02300_ VPWR VGND _04728_ sg13g2_nor2_1
X_24452_ _02325_ _03750_ VPWR VGND _04729_ sg13g2_nor2_1
X_24453_ _03743_ _04728_ _04729_ _03761_ VPWR VGND 
+ _04730_
+ sg13g2_a22oi_1
X_24454_ _02300_ _03763_ VPWR VGND _04731_ sg13g2_nand2b_1
X_24455_ _04237_ _02325_ _04731_ VPWR VGND _04732_ sg13g2_o21ai_1
X_24456_ _03758_ _04732_ _04391_ VPWR VGND _04733_ sg13g2_a21oi_1
X_24457_ _03739_ _04730_ _04733_ VPWR VGND _04734_ sg13g2_a21oi_1
X_24458_ _04727_ _04734_ VPWR VGND _04735_ sg13g2_or2_1
X_24459_ \atbs_core_0.spike_memory_0.n2381_o[12]\ _12085_ VPWR VGND _04736_ sg13g2_nor2_1
X_24460_ \atbs_core_0.spike_memory_0.n2378_o[12]\ _04292_ VPWR VGND _04737_ sg13g2_nor2_1
X_24461_ _03854_ _02246_ VPWR VGND _04738_ sg13g2_nor2_1
X_24462_ _02269_ _03784_ VPWR VGND _04739_ sg13g2_nor2_1
X_24463_ _03842_ _04738_ _04739_ _04051_ VPWR VGND 
+ _04740_
+ sg13g2_a22oi_1
X_24464_ _02246_ _03862_ VPWR VGND _04741_ sg13g2_nand2b_1
X_24465_ _04050_ _02269_ _04741_ VPWR VGND _04742_ sg13g2_o21ai_1
X_24466_ _03757_ _04742_ _03867_ VPWR VGND _04743_ sg13g2_a21oi_1
X_24467_ _03992_ _04740_ _04743_ VPWR VGND _04744_ sg13g2_a21oi_1
X_24468_ _03773_ _04736_ _04737_ _04744_ VPWR VGND 
+ _04745_
+ sg13g2_nor4_1
X_24469_ _07555_ VPWR VGND _04746_ sg13g2_buf_1
X_24470_ \atbs_core_0.spike_memory_0.n2389_o[12]\ _03802_ VPWR VGND _04747_ sg13g2_nor2_1
X_24471_ \atbs_core_0.spike_memory_0.n2386_o[12]\ _04078_ VPWR VGND _04748_ sg13g2_nor2_1
X_24472_ _03988_ _02356_ VPWR VGND _04749_ sg13g2_nor2_1
X_24473_ _02379_ _03850_ VPWR VGND _04750_ sg13g2_nor2_1
X_24474_ _04062_ _04749_ _04750_ _04597_ VPWR VGND 
+ _04751_
+ sg13g2_a22oi_1
X_24475_ _02356_ _03981_ VPWR VGND _04752_ sg13g2_nand2b_1
X_24476_ _03846_ _02379_ _04752_ VPWR VGND _04753_ sg13g2_o21ai_1
X_24477_ _03859_ _04753_ _04068_ VPWR VGND _04754_ sg13g2_a21oi_1
X_24478_ _03839_ _04751_ _04754_ VPWR VGND _04755_ sg13g2_a21oi_1
X_24479_ _04746_ _04747_ _04748_ _04755_ VPWR VGND 
+ _04756_
+ sg13g2_nor4_1
X_24480_ _04745_ _04756_ _04276_ VPWR VGND _04757_ sg13g2_o21ai_1
X_24481_ _04277_ _04735_ _04757_ VPWR VGND _04758_ sg13g2_o21ai_1
X_24482_ _04442_ VPWR VGND _04759_ sg13g2_buf_1
X_24483_ \atbs_core_0.spike_memory_0.n2405_o[12]\ _04759_ VPWR VGND _04760_ sg13g2_nor2_1
X_24484_ \atbs_core_0.spike_memory_0.n2402_o[12]\ _03779_ VPWR VGND _04761_ sg13g2_nor2_1
X_24485_ _04254_ _02584_ VPWR VGND _04762_ sg13g2_nor2_1
X_24486_ _02605_ _03842_ VPWR VGND _04763_ sg13g2_nor2_1
X_24487_ _04108_ _04762_ _04763_ _03983_ VPWR VGND 
+ _04764_
+ sg13g2_a22oi_1
X_24488_ _02584_ _04088_ VPWR VGND _04765_ sg13g2_nand2b_1
X_24489_ _04094_ _02605_ _04765_ VPWR VGND _04766_ sg13g2_o21ai_1
X_24490_ _04010_ _04766_ _03810_ VPWR VGND _04767_ sg13g2_a21oi_1
X_24491_ _04002_ _04764_ _04767_ VPWR VGND _04768_ sg13g2_a21oi_1
X_24492_ _12094_ _04760_ _04761_ _04768_ VPWR VGND 
+ _04769_
+ sg13g2_nor4_1
X_24493_ \atbs_core_0.spike_memory_0.n2401_o[12]\ _12086_ VPWR VGND _04770_ sg13g2_nor2_1
X_24494_ _03778_ VPWR VGND _04771_ sg13g2_buf_1
X_24495_ \atbs_core_0.spike_memory_0.n2398_o[12]\ _04771_ _03780_ VPWR VGND _04772_ sg13g2_o21ai_1
X_24496_ _03787_ _02536_ VPWR VGND _04773_ sg13g2_nor2_1
X_24497_ _02558_ _03785_ VPWR VGND _04774_ sg13g2_nor2_1
X_24498_ _03782_ _04773_ _04774_ _03754_ VPWR VGND 
+ _04775_
+ sg13g2_a22oi_1
X_24499_ _02536_ _03891_ VPWR VGND _04776_ sg13g2_nand2b_1
X_24500_ _03753_ _02558_ _04776_ VPWR VGND _04777_ sg13g2_o21ai_1
X_24501_ _03790_ _04777_ _04294_ VPWR VGND _04778_ sg13g2_a21oi_1
X_24502_ _02700_ _04775_ _04778_ VPWR VGND _04779_ sg13g2_a21oi_1
X_24503_ _04770_ _04772_ _04779_ VPWR VGND _04780_ sg13g2_nor3_1
X_24504_ \atbs_core_0.spike_memory_0.n2397_o[12]\ _03876_ VPWR VGND _04781_ sg13g2_nor2_1
X_24505_ \atbs_core_0.spike_memory_0.n2394_o[12]\ _03835_ VPWR VGND _04782_ sg13g2_nor2_1
X_24506_ _04115_ _02489_ VPWR VGND _04783_ sg13g2_nor2_1
X_24507_ _02510_ _04006_ VPWR VGND _04784_ sg13g2_nor2_1
X_24508_ _04003_ _04783_ _04784_ _03978_ VPWR VGND 
+ _04785_
+ sg13g2_a22oi_1
X_24509_ _02489_ _04110_ VPWR VGND _04786_ sg13g2_nand2b_1
X_24510_ _03760_ _02510_ _04786_ VPWR VGND _04787_ sg13g2_o21ai_1
X_24511_ _04386_ _04787_ _04391_ VPWR VGND _04788_ sg13g2_a21oi_1
X_24512_ _04324_ _04785_ _04788_ VPWR VGND _04789_ sg13g2_a21oi_1
X_24513_ _03727_ _04781_ _04782_ _04789_ VPWR VGND 
+ _04790_
+ sg13g2_nor4_1
X_24514_ _04769_ _04780_ _04790_ VPWR VGND _04791_ sg13g2_or3_1
X_24515_ _03720_ _04758_ _04791_ _03717_ _04335_ VPWR 
+ VGND
+ _04792_ sg13g2_a221oi_1
X_24516_ _12079_ _04725_ _04792_ VPWR VGND _04793_ sg13g2_o21ai_1
X_24517_ _04503_ _04690_ _04793_ VPWR VGND _04794_ sg13g2_nand3_1
X_24518_ _04333_ _04650_ _04794_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[12]\ sg13g2_o21ai_1
X_24519_ _04347_ _02405_ VPWR VGND _04795_ sg13g2_nor2_1
X_24520_ _02424_ _03976_ VPWR VGND _04796_ sg13g2_nor2_1
X_24521_ _04570_ _04795_ _04796_ _04343_ VPWR VGND 
+ _04797_
+ sg13g2_a22oi_1
X_24522_ _02405_ _03788_ VPWR VGND _04798_ sg13g2_nand2b_1
X_24523_ _04347_ _02424_ _04798_ VPWR VGND _04799_ sg13g2_o21ai_1
X_24524_ _03861_ _04799_ _03974_ VPWR VGND _04800_ sg13g2_a21oi_1
X_24525_ _04338_ _04797_ _04800_ VPWR VGND _04801_ sg13g2_a21oi_1
X_24526_ _00150_ _03733_ _03737_ _02459_ _04801_ VPWR 
+ VGND
+ _04802_ sg13g2_a221oi_1
X_24527_ _04357_ _02150_ VPWR VGND _04803_ sg13g2_nor2_1
X_24528_ _02173_ _04359_ VPWR VGND _04804_ sg13g2_nor2_1
X_24529_ _04356_ _04803_ _04804_ _04362_ VPWR VGND 
+ _04805_
+ sg13g2_a22oi_1
X_24530_ _02150_ _03822_ VPWR VGND _04806_ sg13g2_nand2b_1
X_24531_ _04365_ _02173_ _04806_ VPWR VGND _04807_ sg13g2_o21ai_1
X_24532_ _04364_ _04807_ _03740_ VPWR VGND _04808_ sg13g2_a21oi_1
X_24533_ _04355_ _04805_ _04808_ VPWR VGND _04809_ sg13g2_a21oi_1
X_24534_ _00006_ _04353_ _04354_ _02214_ _04809_ VPWR 
+ VGND
+ _04810_ sg13g2_a221oi_1
X_24535_ _00149_ _03969_ VPWR VGND _04811_ sg13g2_nand2_1
X_24536_ \atbs_core_0.spike_memory_0.n2409_o[13]\ _04373_ _04811_ VPWR VGND _04812_ sg13g2_o21ai_1
X_24537_ _04379_ _02632_ VPWR VGND _04813_ sg13g2_nor2_1
X_24538_ _02653_ _04381_ VPWR VGND _04814_ sg13g2_nor2_1
X_24539_ _04511_ _04813_ _04814_ _04384_ VPWR VGND 
+ _04815_
+ sg13g2_a22oi_1
X_24540_ _02632_ _04268_ VPWR VGND _04816_ sg13g2_nand2b_1
X_24541_ _04383_ _02653_ _04816_ VPWR VGND _04817_ sg13g2_o21ai_1
X_24542_ _04517_ _04817_ _04521_ VPWR VGND _04818_ sg13g2_a21oi_1
X_24543_ _04377_ _04815_ _04818_ VPWR VGND _04819_ sg13g2_a21oi_1
X_24544_ _12078_ _04812_ _04819_ VPWR VGND _04820_ sg13g2_nor3_1
X_24545_ _04337_ _04802_ _04810_ _04371_ _04820_ VPWR 
+ VGND
+ _04821_ sg13g2_a221oi_1
X_24546_ \atbs_core_0.spike_memory_0.n2436_q[1210]\ _03776_ VPWR VGND _04822_ sg13g2_nor2_1
X_24547_ \atbs_core_0.spike_memory_0.n2418_o[13]\ _03806_ VPWR VGND _04823_ sg13g2_nor2_1
X_24548_ _03855_ _12646_ VPWR VGND _04824_ sg13g2_nor2_1
X_24549_ _12671_ _03951_ VPWR VGND _04825_ sg13g2_nor2_1
X_24550_ _04047_ _04824_ _04825_ _04052_ VPWR VGND 
+ _04826_
+ sg13g2_a22oi_1
X_24551_ _12646_ _04054_ VPWR VGND _04827_ sg13g2_nand2b_1
X_24552_ _04051_ _12671_ _04827_ VPWR VGND _04828_ sg13g2_o21ai_1
X_24553_ _03955_ _04828_ _03868_ VPWR VGND _04829_ sg13g2_a21oi_1
X_24554_ _03993_ _04826_ _04829_ VPWR VGND _04830_ sg13g2_a21oi_1
X_24555_ _12094_ _04822_ _04823_ _04830_ VPWR VGND 
+ _04831_
+ sg13g2_nor4_1
X_24556_ \atbs_core_0.spike_memory_0.n2417_o[13]\ _04076_ VPWR VGND _04832_ sg13g2_nor2_1
X_24557_ \atbs_core_0.spike_memory_0.n2414_o[13]\ _03835_ _03723_ VPWR VGND _04833_ sg13g2_o21ai_1
X_24558_ _04089_ _12587_ VPWR VGND _04834_ sg13g2_nor2_1
X_24559_ _12611_ _04086_ VPWR VGND _04835_ sg13g2_nor2_1
X_24560_ _04082_ _04834_ _04835_ _04090_ VPWR VGND 
+ _04836_
+ sg13g2_a22oi_1
X_24561_ _12587_ _04094_ VPWR VGND _04837_ sg13g2_nand2b_1
X_24562_ _04413_ _12611_ _04837_ VPWR VGND _04838_ sg13g2_o21ai_1
X_24563_ _04097_ VPWR VGND _04839_ sg13g2_buf_1
X_24564_ _04092_ _04838_ _04839_ VPWR VGND _04840_ sg13g2_a21oi_1
X_24565_ _04081_ _04836_ _04840_ VPWR VGND _04841_ sg13g2_a21oi_1
X_24566_ _04832_ _04833_ _04841_ VPWR VGND _04842_ sg13g2_nor3_1
X_24567_ \atbs_core_0.spike_memory_0.n2413_o[13]\ _03803_ VPWR VGND _04843_ sg13g2_nor2_1
X_24568_ \atbs_core_0.spike_memory_0.n2410_o[13]\ _04102_ VPWR VGND _04844_ sg13g2_nor2_1
X_24569_ _03989_ _12533_ VPWR VGND _04845_ sg13g2_nor2_1
X_24570_ _12555_ _04422_ VPWR VGND _04846_ sg13g2_nor2_1
X_24571_ _04280_ _04845_ _04846_ _04283_ VPWR VGND 
+ _04847_
+ sg13g2_a22oi_1
X_24572_ _12533_ _04425_ VPWR VGND _04848_ sg13g2_nand2b_1
X_24573_ _03847_ _12555_ _04848_ VPWR VGND _04849_ sg13g2_o21ai_1
X_24574_ _03860_ _04849_ _04287_ VPWR VGND _04850_ sg13g2_a21oi_1
X_24575_ _04392_ _04847_ _04850_ VPWR VGND _04851_ sg13g2_a21oi_1
X_24576_ _03800_ _04843_ _04844_ _04851_ VPWR VGND 
+ _04852_
+ sg13g2_nor4_1
X_24577_ _04831_ _04842_ _04852_ VPWR VGND _04853_ sg13g2_nor3_1
X_24578_ \atbs_core_0.spike_memory_0.n2401_o[13]\ _03970_ VPWR VGND _04854_ sg13g2_nand2b_1
X_24579_ \atbs_core_0.spike_memory_0.n2398_o[13]\ _04292_ _04854_ VPWR VGND _04855_ sg13g2_o21ai_1
X_24580_ _04011_ _02537_ VPWR VGND _04856_ sg13g2_nor2_1
X_24581_ _02559_ _04085_ VPWR VGND _04857_ sg13g2_nor2_1
X_24582_ _03750_ _04856_ _04857_ _04413_ VPWR VGND 
+ _04858_
+ sg13g2_a22oi_1
X_24583_ _02537_ _04093_ VPWR VGND _04859_ sg13g2_nand2b_1
X_24584_ _04088_ _02559_ _04859_ VPWR VGND _04860_ sg13g2_o21ai_1
X_24585_ _03986_ _04860_ _04097_ VPWR VGND _04861_ sg13g2_a21oi_1
X_24586_ _03768_ _04858_ _04861_ VPWR VGND _04862_ sg13g2_a21oi_1
X_24587_ _04855_ _04862_ VPWR VGND _04863_ sg13g2_or2_1
X_24588_ \atbs_core_0.spike_memory_0.n2397_o[13]\ _12084_ VPWR VGND _04864_ sg13g2_nor2_1
X_24589_ \atbs_core_0.spike_memory_0.n2394_o[13]\ _03999_ VPWR VGND _04865_ sg13g2_nor2_1
X_24590_ _03890_ _02490_ VPWR VGND _04866_ sg13g2_nor2_1
X_24591_ _02511_ _03741_ VPWR VGND _04867_ sg13g2_nor2_1
X_24592_ _03850_ _04866_ _04867_ _03791_ VPWR VGND 
+ _04868_
+ sg13g2_a22oi_1
X_24593_ _02490_ _02709_ VPWR VGND _04869_ sg13g2_nand2b_1
X_24594_ _03890_ _02511_ _04869_ VPWR VGND _04870_ sg13g2_o21ai_1
X_24595_ _03730_ _04870_ _02698_ VPWR VGND _04871_ sg13g2_a21oi_1
X_24596_ _03867_ _04868_ _04871_ VPWR VGND _04872_ sg13g2_a21oi_1
X_24597_ _03726_ _04864_ _04865_ _04872_ VPWR VGND 
+ _04873_
+ sg13g2_nor4_1
X_24598_ \atbs_core_0.spike_memory_0.n2405_o[13]\ _04442_ VPWR VGND _04874_ sg13g2_nor2_1
X_24599_ \atbs_core_0.spike_memory_0.n2402_o[13]\ _03999_ VPWR VGND _04875_ sg13g2_nor2_1
X_24600_ _04455_ _02585_ VPWR VGND _04876_ sg13g2_nor2_1
X_24601_ _02606_ _03741_ VPWR VGND _04877_ sg13g2_nor2_1
X_24602_ _04085_ _04876_ _04877_ _03915_ VPWR VGND 
+ _04878_
+ sg13g2_a22oi_1
X_24603_ _02585_ _03845_ VPWR VGND _04879_ sg13g2_nand2b_1
X_24604_ _04455_ _02606_ _04879_ VPWR VGND _04880_ sg13g2_o21ai_1
X_24605_ _03730_ _04880_ _03809_ VPWR VGND _04881_ sg13g2_a21oi_1
X_24606_ _04068_ _04878_ _04881_ VPWR VGND _04882_ sg13g2_a21oi_1
X_24607_ _07555_ _04874_ _04875_ _04882_ VPWR VGND 
+ _04883_
+ sg13g2_nor4_1
X_24608_ _04873_ _04883_ _12090_ VPWR VGND _04884_ sg13g2_o21ai_1
X_24609_ _04276_ _04863_ _04884_ VPWR VGND _04885_ sg13g2_o21ai_1
X_24610_ \atbs_core_0.spike_memory_0.n2389_o[13]\ _12085_ VPWR VGND _04886_ sg13g2_nor2_1
X_24611_ \atbs_core_0.spike_memory_0.n2386_o[13]\ _03778_ VPWR VGND _04887_ sg13g2_nor2_1
X_24612_ _03981_ _02357_ VPWR VGND _04888_ sg13g2_nor2_1
X_24613_ _02380_ _03749_ VPWR VGND _04889_ sg13g2_nor2_1
X_24614_ _04107_ _04888_ _04889_ _03863_ VPWR VGND 
+ _04890_
+ sg13g2_a22oi_1
X_24615_ _02357_ _03845_ VPWR VGND _04891_ sg13g2_nand2b_1
X_24616_ _03862_ _02380_ _04891_ VPWR VGND _04892_ sg13g2_o21ai_1
X_24617_ _04009_ _04892_ _03809_ VPWR VGND _04893_ sg13g2_a21oi_1
X_24618_ _04097_ _04890_ _04893_ VPWR VGND _04894_ sg13g2_a21oi_1
X_24619_ _04886_ _04887_ _04894_ VPWR VGND _04895_ sg13g2_nor3_1
X_24620_ \atbs_core_0.spike_memory_0.n2381_o[13]\ _04442_ VPWR VGND _04896_ sg13g2_nor2_1
X_24621_ \atbs_core_0.spike_memory_0.n2378_o[13]\ _03778_ VPWR VGND _04897_ sg13g2_nor2_1
X_24622_ _04093_ _02247_ VPWR VGND _04898_ sg13g2_nor2_1
X_24623_ _02270_ _03749_ VPWR VGND _04899_ sg13g2_nor2_1
X_24624_ _04107_ _04898_ _04899_ _03982_ VPWR VGND 
+ _04900_
+ sg13g2_a22oi_1
X_24625_ _02247_ _03762_ VPWR VGND _04901_ sg13g2_nand2b_1
X_24626_ _03981_ _02270_ _04901_ VPWR VGND _04902_ sg13g2_o21ai_1
X_24627_ _04009_ _04902_ _03767_ VPWR VGND _04903_ sg13g2_a21oi_1
X_24628_ _02699_ _04900_ _04903_ VPWR VGND _04904_ sg13g2_a21oi_1
X_24629_ _03726_ _04896_ _04897_ _04904_ VPWR VGND 
+ _04905_
+ sg13g2_nor4_1
X_24630_ _03727_ _04895_ _04905_ VPWR VGND _04906_ sg13g2_a21oi_1
X_24631_ _03745_ _02302_ VPWR VGND _04907_ sg13g2_nor2_1
X_24632_ _02326_ _03784_ VPWR VGND _04908_ sg13g2_nor2_1
X_24633_ _03742_ _04907_ _04908_ _03787_ VPWR VGND 
+ _04909_
+ sg13g2_a22oi_1
X_24634_ _02302_ _03890_ VPWR VGND _04910_ sg13g2_nand2b_1
X_24635_ _03745_ _02326_ _04910_ VPWR VGND _04911_ sg13g2_o21ai_1
X_24636_ _03757_ _04911_ _03767_ VPWR VGND _04912_ sg13g2_a21oi_1
X_24637_ _03738_ _04909_ _04912_ VPWR VGND _04913_ sg13g2_a21oi_1
X_24638_ \atbs_core_0.spike_memory_0.n2385_o[13]\ _12085_ _07552_ VPWR VGND _04914_ sg13g2_o21ai_1
X_24639_ _07555_ _04913_ _04914_ VPWR VGND _04915_ sg13g2_nor3_1
X_24640_ \atbs_core_0.spike_memory_0.n2382_o[13]\ _04230_ _04915_ VPWR VGND _04916_ sg13g2_o21ai_1
X_24641_ _03966_ _04906_ _04916_ VPWR VGND _04917_ sg13g2_o21ai_1
X_24642_ _07541_ _04885_ _04917_ _03720_ VPWR VGND 
+ _04918_
+ sg13g2_a22oi_1
X_24643_ _12079_ _04853_ _04918_ VPWR VGND _04919_ sg13g2_o21ai_1
X_24644_ _04336_ _04919_ VPWR VGND _04920_ sg13g2_nor2_1
X_24645_ _04336_ _04821_ _04920_ VPWR VGND _04921_ sg13g2_a21oi_1
X_24646_ \atbs_core_0.spike_memory_0.n2361_o[13]\ _04506_ VPWR VGND _04922_ sg13g2_nor2_1
X_24647_ \atbs_core_0.spike_memory_0.n2358_o[13]\ _04508_ VPWR VGND _04923_ sg13g2_nor2_1
X_24648_ _04513_ _02142_ VPWR VGND _04924_ sg13g2_nor2_1
X_24649_ _02334_ _04381_ VPWR VGND _04925_ sg13g2_nor2_1
X_24650_ _04511_ _04924_ _04925_ _04384_ VPWR VGND 
+ _04926_
+ sg13g2_a22oi_1
X_24651_ _02142_ _04518_ VPWR VGND _04927_ sg13g2_nand2b_1
X_24652_ _04383_ _02334_ _04927_ VPWR VGND _04928_ sg13g2_o21ai_1
X_24653_ _04517_ _04928_ _04521_ VPWR VGND _04929_ sg13g2_a21oi_1
X_24654_ _04377_ _04926_ _04929_ VPWR VGND _04930_ sg13g2_a21oi_1
X_24655_ _04505_ _04922_ _04923_ _04930_ VPWR VGND 
+ _04931_
+ sg13g2_nor4_1
X_24656_ \atbs_core_0.spike_memory_0.n2369_o[13]\ _04525_ VPWR VGND _04932_ sg13g2_nor2_1
X_24657_ \atbs_core_0.spike_memory_0.n2366_o[13]\ _04528_ VPWR VGND _04933_ sg13g2_nor2_1
X_24658_ _03887_ _02040_ VPWR VGND _04934_ sg13g2_nor2_1
X_24659_ _02062_ _04533_ VPWR VGND _04935_ sg13g2_nor2_1
X_24660_ _04531_ _04934_ _04935_ _04536_ VPWR VGND 
+ _04936_
+ sg13g2_a22oi_1
X_24661_ _02040_ _04559_ VPWR VGND _04937_ sg13g2_nand2b_1
X_24662_ _04539_ _02062_ _04937_ VPWR VGND _04938_ sg13g2_o21ai_1
X_24663_ _04538_ _04938_ _04542_ VPWR VGND _04939_ sg13g2_a21oi_1
X_24664_ _04530_ _04936_ _04939_ VPWR VGND _04940_ sg13g2_a21oi_1
X_24665_ _04604_ _04932_ _04933_ _04940_ VPWR VGND 
+ _04941_
+ sg13g2_nor4_1
X_24666_ _04504_ _04931_ _04941_ VPWR VGND _04942_ sg13g2_nor3_1
X_24667_ \atbs_core_0.spike_memory_0.n2365_o[13]\ _04525_ VPWR VGND _04943_ sg13g2_nor2_1
X_24668_ \atbs_core_0.spike_memory_0.n2362_o[13]\ _04549_ VPWR VGND _04944_ sg13g2_nor2_1
X_24669_ _04553_ _12580_ VPWR VGND _04945_ sg13g2_nor2_1
X_24670_ _02013_ _04555_ VPWR VGND _04946_ sg13g2_nor2_1
X_24671_ _04378_ _04945_ _04946_ _04557_ VPWR VGND 
+ _04947_
+ sg13g2_a22oi_1
X_24672_ _12580_ _04559_ VPWR VGND _04948_ sg13g2_nand2b_1
X_24673_ _03755_ _02013_ _04948_ VPWR VGND _04949_ sg13g2_o21ai_1
X_24674_ _04388_ _04949_ _04562_ VPWR VGND _04950_ sg13g2_a21oi_1
X_24675_ _04551_ _04947_ _04950_ VPWR VGND _04951_ sg13g2_a21oi_1
X_24676_ _03729_ _04943_ _04944_ _04951_ VPWR VGND 
+ _04952_
+ sg13g2_nor4_1
X_24677_ \atbs_core_0.spike_memory_0.n2373_o[13]\ _12088_ VPWR VGND _04953_ sg13g2_nor2_1
X_24678_ \atbs_core_0.spike_memory_0.n2370_o[13]\ _04528_ VPWR VGND _04954_ sg13g2_nor2_1
X_24679_ _03934_ _02095_ VPWR VGND _04955_ sg13g2_nor2_1
X_24680_ _02117_ _04570_ VPWR VGND _04956_ sg13g2_nor2_1
X_24681_ _04568_ _04955_ _04956_ _02714_ VPWR VGND 
+ _04957_
+ sg13g2_a22oi_1
X_24682_ _02095_ _04361_ VPWR VGND _04958_ sg13g2_nand2b_1
X_24683_ _04574_ _02117_ _04958_ VPWR VGND _04959_ sg13g2_o21ai_1
X_24684_ _04573_ _04959_ _04338_ VPWR VGND _04960_ sg13g2_a21oi_1
X_24685_ _02702_ _04957_ _04960_ VPWR VGND _04961_ sg13g2_a21oi_1
X_24686_ _04126_ _04953_ _04954_ _04961_ VPWR VGND 
+ _04962_
+ sg13g2_nor4_1
X_24687_ _04547_ _04952_ _04962_ VPWR VGND _04963_ sg13g2_nor3_1
X_24688_ _04503_ _04942_ _04963_ VPWR VGND _04964_ sg13g2_nor3_1
X_24689_ _04333_ _04921_ _04964_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[13]\ sg13g2_a21o_1
X_24690_ \atbs_core_0.spike_memory_0.n2365_o[14]\ _04582_ VPWR VGND _04965_ sg13g2_nor2_1
X_24691_ \atbs_core_0.spike_memory_0.n2362_o[14]\ _04584_ VPWR VGND _04966_ sg13g2_nor2_1
X_24692_ _04590_ _12592_ VPWR VGND _04967_ sg13g2_nor2_1
X_24693_ _02015_ _04150_ VPWR VGND _04968_ sg13g2_nor2_1
X_24694_ _04588_ _04967_ _04968_ _04594_ VPWR VGND 
+ _04969_
+ sg13g2_a22oi_1
X_24695_ _12592_ _04598_ VPWR VGND _04970_ sg13g2_nand2b_1
X_24696_ _04593_ _02015_ _04970_ VPWR VGND _04971_ sg13g2_o21ai_1
X_24697_ _04596_ _04971_ _02701_ VPWR VGND _04972_ sg13g2_a21oi_1
X_24698_ _04586_ _04969_ _04972_ VPWR VGND _04973_ sg13g2_a21oi_1
X_24699_ _04505_ _04965_ _04966_ _04973_ VPWR VGND 
+ _04974_
+ sg13g2_nor4_1
X_24700_ \atbs_core_0.spike_memory_0.n2373_o[14]\ _04373_ VPWR VGND _04975_ sg13g2_nor2_1
X_24701_ \atbs_core_0.spike_memory_0.n2370_o[14]\ _04606_ VPWR VGND _04976_ sg13g2_nor2_1
X_24702_ _04610_ _02096_ VPWR VGND _04977_ sg13g2_nor2_1
X_24703_ _02119_ _03814_ VPWR VGND _04978_ sg13g2_nor2_1
X_24704_ _04609_ _04977_ _04978_ _04613_ VPWR VGND 
+ _04979_
+ sg13g2_a22oi_1
X_24705_ _02096_ _04283_ VPWR VGND _04980_ sg13g2_nand2b_1
X_24706_ _04616_ _02119_ _04980_ VPWR VGND _04981_ sg13g2_o21ai_1
X_24707_ _04615_ _04981_ _03948_ VPWR VGND _04982_ sg13g2_a21oi_1
X_24708_ _04608_ _04979_ _04982_ VPWR VGND _04983_ sg13g2_a21oi_1
X_24709_ _04604_ _04975_ _04976_ _04983_ VPWR VGND 
+ _04984_
+ sg13g2_nor4_1
X_24710_ _04974_ _04984_ _04504_ VPWR VGND _04985_ sg13g2_o21ai_1
X_24711_ \atbs_core_0.spike_memory_0.n2361_o[14]\ _04623_ VPWR VGND _04986_ sg13g2_nor2_1
X_24712_ \atbs_core_0.spike_memory_0.n2358_o[14]\ _04584_ VPWR VGND _04987_ sg13g2_nor2_1
X_24713_ _04593_ _02154_ VPWR VGND _04988_ sg13g2_nor2_1
X_24714_ _02336_ _04628_ VPWR VGND _04989_ sg13g2_nor2_1
X_24715_ _04588_ _04988_ _04989_ _04630_ VPWR VGND 
+ _04990_
+ sg13g2_a22oi_1
X_24716_ _02154_ _04052_ VPWR VGND _04991_ sg13g2_nand2b_1
X_24717_ _04632_ _02336_ _04991_ VPWR VGND _04992_ sg13g2_o21ai_1
X_24718_ _04596_ _04992_ _04635_ VPWR VGND _04993_ sg13g2_a21oi_1
X_24719_ _04626_ _04990_ _04993_ VPWR VGND _04994_ sg13g2_a21oi_1
X_24720_ _03872_ _04986_ _04987_ _04994_ VPWR VGND 
+ _04995_
+ sg13g2_nor4_1
X_24721_ \atbs_core_0.spike_memory_0.n2369_o[14]\ _04582_ VPWR VGND _04996_ sg13g2_nor2_1
X_24722_ \atbs_core_0.spike_memory_0.n2366_o[14]\ _04606_ VPWR VGND _04997_ sg13g2_nor2_1
X_24723_ _04616_ _02041_ VPWR VGND _04998_ sg13g2_nor2_1
X_24724_ _02063_ _04035_ VPWR VGND _04999_ sg13g2_nor2_1
X_24725_ _04609_ _04998_ _04999_ _04594_ VPWR VGND 
+ _05000_
+ sg13g2_a22oi_1
X_24726_ _02041_ _03848_ VPWR VGND _05001_ sg13g2_nand2b_1
X_24727_ _04590_ _02063_ _05001_ VPWR VGND _05002_ sg13g2_o21ai_1
X_24728_ _04615_ _05002_ _04149_ VPWR VGND _05003_ sg13g2_a21oi_1
X_24729_ _04586_ _05000_ _05003_ VPWR VGND _05004_ sg13g2_a21oi_1
X_24730_ _04219_ _04996_ _04997_ _05004_ VPWR VGND 
+ _05005_
+ sg13g2_nor4_1
X_24731_ _04995_ _05005_ _04547_ VPWR VGND _05006_ sg13g2_o21ai_1
X_24732_ _04985_ _05006_ VPWR VGND _05007_ sg13g2_and2_1
X_24733_ _04651_ _02406_ VPWR VGND _05008_ sg13g2_nor2_1
X_24734_ _02425_ _04510_ VPWR VGND _05009_ sg13g2_nor2_1
X_24735_ _04356_ _05008_ _05009_ _04680_ VPWR VGND 
+ _05010_
+ sg13g2_a22oi_1
X_24736_ _02406_ _03882_ VPWR VGND _05011_ sg13g2_nand2b_1
X_24737_ _04320_ _02425_ _05011_ VPWR VGND _05012_ sg13g2_o21ai_1
X_24738_ _04364_ _05012_ _04376_ VPWR VGND _05013_ sg13g2_a21oi_1
X_24739_ _04677_ _05010_ _05013_ VPWR VGND _05014_ sg13g2_a21oi_1
X_24740_ _00008_ _04675_ _04676_ _02461_ _05014_ VPWR 
+ VGND
+ _05015_ sg13g2_a221oi_1
X_24741_ _04632_ _02633_ VPWR VGND _05016_ sg13g2_nor2_1
X_24742_ _02655_ _04628_ VPWR VGND _05017_ sg13g2_nor2_1
X_24743_ _04662_ _05016_ _05017_ _04630_ VPWR VGND 
+ _05018_
+ sg13g2_a22oi_1
X_24744_ _02633_ _03957_ VPWR VGND _05019_ sg13g2_nand2b_1
X_24745_ _04365_ _02655_ _05019_ VPWR VGND _05020_ sg13g2_o21ai_1
X_24746_ _04666_ _05020_ _03880_ VPWR VGND _05021_ sg13g2_a21oi_1
X_24747_ _04626_ _05018_ _05021_ VPWR VGND _05022_ sg13g2_a21oi_1
X_24748_ _00007_ _04660_ _04661_ _02685_ _05022_ VPWR 
+ VGND
+ _05023_ sg13g2_a221oi_1
X_24749_ _04337_ _05015_ _05023_ _04673_ VPWR VGND 
+ _05024_
+ sg13g2_a22oi_1
X_24750_ _04651_ _02151_ VPWR VGND _05025_ sg13g2_nor2_1
X_24751_ _02174_ _04510_ VPWR VGND _05026_ sg13g2_nor2_1
X_24752_ _04339_ _05025_ _05026_ _04680_ VPWR VGND 
+ _05027_
+ sg13g2_a22oi_1
X_24753_ _02151_ _04552_ VPWR VGND _05028_ sg13g2_nand2b_1
X_24754_ _04340_ _02174_ _05028_ VPWR VGND _05029_ sg13g2_o21ai_1
X_24755_ _04345_ _05029_ _04684_ VPWR VGND _05030_ sg13g2_a21oi_1
X_24756_ _04677_ _05027_ _05030_ VPWR VGND _05031_ sg13g2_a21oi_1
X_24757_ _00009_ _04675_ _04676_ _02216_ _05031_ VPWR 
+ VGND
+ _05032_ sg13g2_a221oi_1
X_24758_ _04371_ _05032_ _04688_ VPWR VGND _05033_ sg13g2_a21oi_1
X_24759_ _05024_ _05033_ VPWR VGND _05034_ sg13g2_nand2_1
X_24760_ \atbs_core_0.spike_memory_0.n2413_o[14]\ _03901_ VPWR VGND _05035_ sg13g2_nor2_1
X_24761_ \atbs_core_0.spike_memory_0.n2410_o[14]\ _03807_ VPWR VGND _05036_ sg13g2_nor2_1
X_24762_ _03816_ _12534_ VPWR VGND _05037_ sg13g2_nor2_1
X_24763_ _12557_ _03819_ VPWR VGND _05038_ sg13g2_nor2_1
X_24764_ _04035_ _05037_ _05038_ _03823_ VPWR VGND 
+ _05039_
+ sg13g2_a22oi_1
X_24765_ _12534_ _03916_ VPWR VGND _05040_ sg13g2_nand2b_1
X_24766_ _03930_ _12557_ _05040_ VPWR VGND _05041_ sg13g2_o21ai_1
X_24767_ _03825_ _05041_ _04142_ VPWR VGND _05042_ sg13g2_a21oi_1
X_24768_ _03812_ _05039_ _05042_ VPWR VGND _05043_ sg13g2_a21oi_1
X_24769_ _04074_ _05035_ _05036_ _05043_ VPWR VGND 
+ _05044_
+ sg13g2_nor4_1
X_24770_ \atbs_core_0.spike_memory_0.n2417_o[14]\ _04623_ VPWR VGND _05045_ sg13g2_nor2_1
X_24771_ \atbs_core_0.spike_memory_0.n2414_o[14]\ _04702_ _03966_ VPWR VGND _05046_ sg13g2_o21ai_1
X_24772_ _04704_ _12589_ VPWR VGND _05047_ sg13g2_nor2_1
X_24773_ _12612_ _04587_ VPWR VGND _05048_ sg13g2_nor2_1
X_24774_ _04381_ _05047_ _05048_ _04343_ VPWR VGND 
+ _05049_
+ sg13g2_a22oi_1
X_24775_ _12589_ _04589_ VPWR VGND _05050_ sg13g2_nand2b_1
X_24776_ _04708_ _12612_ _05050_ VPWR VGND _05051_ sg13g2_o21ai_1
X_24777_ _03861_ _05051_ _03869_ VPWR VGND _05052_ sg13g2_a21oi_1
X_24778_ _04393_ _05049_ _05052_ VPWR VGND _05053_ sg13g2_a21oi_1
X_24779_ _05045_ _05046_ _05053_ VPWR VGND _05054_ sg13g2_nor3_1
X_24780_ \atbs_core_0.spike_memory_0.n2436_q[1211]\ _03804_ VPWR VGND _05055_ sg13g2_nor2_1
X_24781_ \atbs_core_0.spike_memory_0.n2418_o[14]\ _03946_ VPWR VGND _05056_ sg13g2_nor2_1
X_24782_ _03848_ _12647_ VPWR VGND _05057_ sg13g2_nor2_1
X_24783_ _12672_ _03852_ VPWR VGND _05058_ sg13g2_nor2_1
X_24784_ _04716_ _05057_ _05058_ _03857_ VPWR VGND 
+ _05059_
+ sg13g2_a22oi_1
X_24785_ _12647_ _03864_ VPWR VGND _05060_ sg13g2_nand2b_1
X_24786_ _04598_ _12672_ _05060_ VPWR VGND _05061_ sg13g2_o21ai_1
X_24787_ _03956_ _05061_ _04317_ VPWR VGND _05062_ sg13g2_a21oi_1
X_24788_ _03841_ _05059_ _05062_ VPWR VGND _05063_ sg13g2_a21oi_1
X_24789_ _12095_ _05055_ _05056_ _05063_ VPWR VGND 
+ _05064_
+ sg13g2_nor4_1
X_24790_ _05044_ _05054_ _05064_ VPWR VGND _05065_ sg13g2_nor3_1
X_24791_ \atbs_core_0.spike_memory_0.n2385_o[14]\ _03970_ VPWR VGND _05066_ sg13g2_nand2b_1
X_24792_ \atbs_core_0.spike_memory_0.n2382_o[14]\ _04771_ _05066_ VPWR VGND _05067_ sg13g2_o21ai_1
X_24793_ _03746_ _02303_ VPWR VGND _05068_ sg13g2_nor2_1
X_24794_ _02327_ _03750_ VPWR VGND _05069_ sg13g2_nor2_1
X_24795_ _03743_ _05068_ _05069_ _03761_ VPWR VGND 
+ _05070_
+ sg13g2_a22oi_1
X_24796_ _02303_ _04110_ VPWR VGND _05071_ sg13g2_nand2b_1
X_24797_ _04237_ _02327_ _05071_ VPWR VGND _05072_ sg13g2_o21ai_1
X_24798_ _04386_ _05072_ _04391_ VPWR VGND _05073_ sg13g2_a21oi_1
X_24799_ _04324_ _05070_ _05073_ VPWR VGND _05074_ sg13g2_a21oi_1
X_24800_ _05067_ _05074_ VPWR VGND _05075_ sg13g2_or2_1
X_24801_ \atbs_core_0.spike_memory_0.n2381_o[14]\ _12085_ VPWR VGND _05076_ sg13g2_nor2_1
X_24802_ \atbs_core_0.spike_memory_0.n2378_o[14]\ _04292_ VPWR VGND _05077_ sg13g2_nor2_1
X_24803_ _03854_ _02248_ VPWR VGND _05078_ sg13g2_nor2_1
X_24804_ _02271_ _03784_ VPWR VGND _05079_ sg13g2_nor2_1
X_24805_ _03842_ _05078_ _05079_ _04051_ VPWR VGND 
+ _05080_
+ sg13g2_a22oi_1
X_24806_ _02248_ _04455_ VPWR VGND _05081_ sg13g2_nand2b_1
X_24807_ _04050_ _02271_ _05081_ VPWR VGND _05082_ sg13g2_o21ai_1
X_24808_ _03757_ _05082_ _03867_ VPWR VGND _05083_ sg13g2_a21oi_1
X_24809_ _03992_ _05080_ _05083_ VPWR VGND _05084_ sg13g2_a21oi_1
X_24810_ _03773_ _05076_ _05077_ _05084_ VPWR VGND 
+ _05085_
+ sg13g2_nor4_1
X_24811_ \atbs_core_0.spike_memory_0.n2389_o[14]\ _03802_ VPWR VGND _05086_ sg13g2_nor2_1
X_24812_ \atbs_core_0.spike_memory_0.n2386_o[14]\ _04078_ VPWR VGND _05087_ sg13g2_nor2_1
X_24813_ _03988_ _02358_ VPWR VGND _05088_ sg13g2_nor2_1
X_24814_ _02381_ _03850_ VPWR VGND _05089_ sg13g2_nor2_1
X_24815_ _04062_ _05088_ _05089_ _04597_ VPWR VGND 
+ _05090_
+ sg13g2_a22oi_1
X_24816_ _02358_ _03981_ VPWR VGND _05091_ sg13g2_nand2b_1
X_24817_ _03846_ _02381_ _05091_ VPWR VGND _05092_ sg13g2_o21ai_1
X_24818_ _03859_ _05092_ _04068_ VPWR VGND _05093_ sg13g2_a21oi_1
X_24819_ _03839_ _05090_ _05093_ VPWR VGND _05094_ sg13g2_a21oi_1
X_24820_ _04746_ _05086_ _05087_ _05094_ VPWR VGND 
+ _05095_
+ sg13g2_nor4_1
X_24821_ _05085_ _05095_ _04276_ VPWR VGND _05096_ sg13g2_o21ai_1
X_24822_ _04277_ _05075_ _05096_ VPWR VGND _05097_ sg13g2_o21ai_1
X_24823_ \atbs_core_0.spike_memory_0.n2405_o[14]\ _04759_ VPWR VGND _05098_ sg13g2_nor2_1
X_24824_ \atbs_core_0.spike_memory_0.n2402_o[14]\ _03779_ VPWR VGND _05099_ sg13g2_nor2_1
X_24825_ _04254_ _02586_ VPWR VGND _05100_ sg13g2_nor2_1
X_24826_ _02607_ _03842_ VPWR VGND _05101_ sg13g2_nor2_1
X_24827_ _04108_ _05100_ _05101_ _03983_ VPWR VGND 
+ _05102_
+ sg13g2_a22oi_1
X_24828_ _02586_ _04088_ VPWR VGND _05103_ sg13g2_nand2b_1
X_24829_ _04094_ _02607_ _05103_ VPWR VGND _05104_ sg13g2_o21ai_1
X_24830_ _04010_ _05104_ _03810_ VPWR VGND _05105_ sg13g2_a21oi_1
X_24831_ _04118_ _05102_ _05105_ VPWR VGND _05106_ sg13g2_a21oi_1
X_24832_ _12093_ _05098_ _05099_ _05106_ VPWR VGND 
+ _05107_
+ sg13g2_nor4_1
X_24833_ \atbs_core_0.spike_memory_0.n2401_o[14]\ _12086_ VPWR VGND _05108_ sg13g2_nor2_1
X_24834_ \atbs_core_0.spike_memory_0.n2398_o[14]\ _04771_ _03780_ VPWR VGND _05109_ sg13g2_o21ai_1
X_24835_ _03787_ _02539_ VPWR VGND _05110_ sg13g2_nor2_1
X_24836_ _02560_ _03785_ VPWR VGND _05111_ sg13g2_nor2_1
X_24837_ _03782_ _05110_ _05111_ _03754_ VPWR VGND 
+ _05112_
+ sg13g2_a22oi_1
X_24838_ _02539_ _03891_ VPWR VGND _05113_ sg13g2_nand2b_1
X_24839_ _03753_ _02560_ _05113_ VPWR VGND _05114_ sg13g2_o21ai_1
X_24840_ _03758_ _05114_ _04294_ VPWR VGND _05115_ sg13g2_a21oi_1
X_24841_ _03739_ _05112_ _05115_ VPWR VGND _05116_ sg13g2_a21oi_1
X_24842_ _05108_ _05109_ _05116_ VPWR VGND _05117_ sg13g2_nor3_1
X_24843_ \atbs_core_0.spike_memory_0.n2397_o[14]\ _03876_ VPWR VGND _05118_ sg13g2_nor2_1
X_24844_ \atbs_core_0.spike_memory_0.n2394_o[14]\ _03835_ VPWR VGND _05119_ sg13g2_nor2_1
X_24845_ _04115_ _02491_ VPWR VGND _05120_ sg13g2_nor2_1
X_24846_ _02512_ _04006_ VPWR VGND _05121_ sg13g2_nor2_1
X_24847_ _04003_ _05120_ _05121_ _03978_ VPWR VGND 
+ _05122_
+ sg13g2_a22oi_1
X_24848_ _02491_ _04110_ VPWR VGND _05123_ sg13g2_nand2b_1
X_24849_ _03760_ _02512_ _05123_ VPWR VGND _05124_ sg13g2_o21ai_1
X_24850_ _04386_ _05124_ _04391_ VPWR VGND _05125_ sg13g2_a21oi_1
X_24851_ _04324_ _05122_ _05125_ VPWR VGND _05126_ sg13g2_a21oi_1
X_24852_ _03727_ _05118_ _05119_ _05126_ VPWR VGND 
+ _05127_
+ sg13g2_nor4_1
X_24853_ _05107_ _05117_ _05127_ VPWR VGND _05128_ sg13g2_or3_1
X_24854_ _03720_ _05097_ _05128_ _03717_ _04335_ VPWR 
+ VGND
+ _05129_ sg13g2_a221oi_1
X_24855_ _12079_ _05065_ _05129_ VPWR VGND _05130_ sg13g2_o21ai_1
X_24856_ _04503_ _05034_ _05130_ VPWR VGND _05131_ sg13g2_nand3_1
X_24857_ _04333_ _05007_ _05131_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[14]\ sg13g2_o21ai_1
X_24858_ \atbs_core_0.spike_memory_0.n2365_o[15]\ _04582_ VPWR VGND _05132_ sg13g2_nor2_1
X_24859_ \atbs_core_0.spike_memory_0.n2362_o[15]\ _04584_ VPWR VGND _05133_ sg13g2_nor2_1
X_24860_ _04590_ _12604_ VPWR VGND _05134_ sg13g2_nor2_1
X_24861_ _02016_ _04150_ VPWR VGND _05135_ sg13g2_nor2_1
X_24862_ _04588_ _05134_ _05135_ _04594_ VPWR VGND 
+ _05136_
+ sg13g2_a22oi_1
X_24863_ _12604_ _04598_ VPWR VGND _05137_ sg13g2_nand2b_1
X_24864_ _04593_ _02016_ _05137_ VPWR VGND _05138_ sg13g2_o21ai_1
X_24865_ _04596_ _05138_ _04635_ VPWR VGND _05139_ sg13g2_a21oi_1
X_24866_ _04586_ _05136_ _05139_ VPWR VGND _05140_ sg13g2_a21oi_1
X_24867_ _03872_ _05132_ _05133_ _05140_ VPWR VGND 
+ _05141_
+ sg13g2_nor4_1
X_24868_ \atbs_core_0.spike_memory_0.n2373_o[15]\ _04373_ VPWR VGND _05142_ sg13g2_nor2_1
X_24869_ \atbs_core_0.spike_memory_0.n2370_o[15]\ _04606_ VPWR VGND _05143_ sg13g2_nor2_1
X_24870_ _04610_ _02097_ VPWR VGND _05144_ sg13g2_nor2_1
X_24871_ _02121_ _03814_ VPWR VGND _05145_ sg13g2_nor2_1
X_24872_ _04609_ _05144_ _05145_ _04613_ VPWR VGND 
+ _05146_
+ sg13g2_a22oi_1
X_24873_ _02097_ _04283_ VPWR VGND _05147_ sg13g2_nand2b_1
X_24874_ _04616_ _02121_ _05147_ VPWR VGND _05148_ sg13g2_o21ai_1
X_24875_ _04615_ _05148_ _03812_ VPWR VGND _05149_ sg13g2_a21oi_1
X_24876_ _04608_ _05146_ _05149_ VPWR VGND _05150_ sg13g2_a21oi_1
X_24877_ _04219_ _05142_ _05143_ _05150_ VPWR VGND 
+ _05151_
+ sg13g2_nor4_1
X_24878_ _05141_ _05151_ _04504_ VPWR VGND _05152_ sg13g2_o21ai_1
X_24879_ \atbs_core_0.spike_memory_0.n2361_o[15]\ _04623_ VPWR VGND _05153_ sg13g2_nor2_1
X_24880_ \atbs_core_0.spike_memory_0.n2358_o[15]\ _04584_ VPWR VGND _05154_ sg13g2_nor2_1
X_24881_ _04593_ _02166_ VPWR VGND _05155_ sg13g2_nor2_1
X_24882_ _02338_ _04628_ VPWR VGND _05156_ sg13g2_nor2_1
X_24883_ _04662_ _05155_ _05156_ _04630_ VPWR VGND 
+ _05157_
+ sg13g2_a22oi_1
X_24884_ _02166_ _04052_ VPWR VGND _05158_ sg13g2_nand2b_1
X_24885_ _04632_ _02338_ _05158_ VPWR VGND _05159_ sg13g2_o21ai_1
X_24886_ _04666_ _05159_ _04635_ VPWR VGND _05160_ sg13g2_a21oi_1
X_24887_ _04626_ _05157_ _05160_ VPWR VGND _05161_ sg13g2_a21oi_1
X_24888_ _03872_ _05153_ _05154_ _05161_ VPWR VGND 
+ _05162_
+ sg13g2_nor4_1
X_24889_ \atbs_core_0.spike_memory_0.n2369_o[15]\ _04582_ VPWR VGND _05163_ sg13g2_nor2_1
X_24890_ \atbs_core_0.spike_memory_0.n2366_o[15]\ _04606_ VPWR VGND _05164_ sg13g2_nor2_1
X_24891_ _04616_ _02042_ VPWR VGND _05165_ sg13g2_nor2_1
X_24892_ _02064_ _04035_ VPWR VGND _05166_ sg13g2_nor2_1
X_24893_ _04588_ _05165_ _05166_ _04594_ VPWR VGND 
+ _05167_
+ sg13g2_a22oi_1
X_24894_ _02042_ _03856_ VPWR VGND _05168_ sg13g2_nand2b_1
X_24895_ _04590_ _02064_ _05168_ VPWR VGND _05169_ sg13g2_o21ai_1
X_24896_ _04596_ _05169_ _04149_ VPWR VGND _05170_ sg13g2_a21oi_1
X_24897_ _04586_ _05167_ _05170_ VPWR VGND _05171_ sg13g2_a21oi_1
X_24898_ _04219_ _05163_ _05164_ _05171_ VPWR VGND 
+ _05172_
+ sg13g2_nor4_1
X_24899_ _05162_ _05172_ _03725_ VPWR VGND _05173_ sg13g2_o21ai_1
X_24900_ _05152_ _05173_ VPWR VGND _05174_ sg13g2_and2_1
X_24901_ _04651_ _02407_ VPWR VGND _05175_ sg13g2_nor2_1
X_24902_ _02426_ _04510_ VPWR VGND _05176_ sg13g2_nor2_1
X_24903_ _04356_ _05175_ _05176_ _04680_ VPWR VGND 
+ _05177_
+ sg13g2_a22oi_1
X_24904_ _02407_ _04552_ VPWR VGND _05178_ sg13g2_nand2b_1
X_24905_ _04320_ _02426_ _05178_ VPWR VGND _05179_ sg13g2_o21ai_1
X_24906_ _04364_ _05179_ _04376_ VPWR VGND _05180_ sg13g2_a21oi_1
X_24907_ _04677_ _05177_ _05180_ VPWR VGND _05181_ sg13g2_a21oi_1
X_24908_ _00011_ _04675_ _04676_ _02463_ _05181_ VPWR 
+ VGND
+ _05182_ sg13g2_a221oi_1
X_24909_ _04632_ _02635_ VPWR VGND _05183_ sg13g2_nor2_1
X_24910_ _02656_ _03881_ VPWR VGND _05184_ sg13g2_nor2_1
X_24911_ _04662_ _05183_ _05184_ _04630_ VPWR VGND 
+ _05185_
+ sg13g2_a22oi_1
X_24912_ _02635_ _03957_ VPWR VGND _05186_ sg13g2_nand2b_1
X_24913_ _04365_ _02656_ _05186_ VPWR VGND _05187_ sg13g2_o21ai_1
X_24914_ _04666_ _05187_ _03880_ VPWR VGND _05188_ sg13g2_a21oi_1
X_24915_ _04626_ _05185_ _05188_ VPWR VGND _05189_ sg13g2_a21oi_1
X_24916_ _00010_ _04660_ _04661_ _02687_ _05189_ VPWR 
+ VGND
+ _05190_ sg13g2_a221oi_1
X_24917_ _04337_ _05182_ _05190_ _04673_ VPWR VGND 
+ _05191_
+ sg13g2_a22oi_1
X_24918_ _04651_ _02152_ VPWR VGND _05192_ sg13g2_nor2_1
X_24919_ _02175_ _03976_ VPWR VGND _05193_ sg13g2_nor2_1
X_24920_ _04339_ _05192_ _05193_ _04680_ VPWR VGND 
+ _05194_
+ sg13g2_a22oi_1
X_24921_ _02152_ _04552_ VPWR VGND _05195_ sg13g2_nand2b_1
X_24922_ _04340_ _02175_ _05195_ VPWR VGND _05196_ sg13g2_o21ai_1
X_24923_ _04345_ _05196_ _04684_ VPWR VGND _05197_ sg13g2_a21oi_1
X_24924_ _04677_ _05194_ _05197_ VPWR VGND _05198_ sg13g2_a21oi_1
X_24925_ _00012_ _04675_ _04676_ _02219_ _05198_ VPWR 
+ VGND
+ _05199_ sg13g2_a221oi_1
X_24926_ _04371_ _05199_ _04688_ VPWR VGND _05200_ sg13g2_a21oi_1
X_24927_ _05191_ _05200_ VPWR VGND _05201_ sg13g2_nand2_1
X_24928_ \atbs_core_0.spike_memory_0.n2413_o[15]\ _03901_ VPWR VGND _05202_ sg13g2_nor2_1
X_24929_ \atbs_core_0.spike_memory_0.n2410_o[15]\ _03903_ VPWR VGND _05203_ sg13g2_nor2_1
X_24930_ _03816_ _12535_ VPWR VGND _05204_ sg13g2_nor2_1
X_24931_ _12558_ _03819_ VPWR VGND _05205_ sg13g2_nor2_1
X_24932_ _04035_ _05204_ _05205_ _03911_ VPWR VGND 
+ _05206_
+ sg13g2_a22oi_1
X_24933_ _12535_ _03916_ VPWR VGND _05207_ sg13g2_nand2b_1
X_24934_ _03930_ _12558_ _05207_ VPWR VGND _05208_ sg13g2_o21ai_1
X_24935_ _03825_ _05208_ _04142_ VPWR VGND _05209_ sg13g2_a21oi_1
X_24936_ _03812_ _05206_ _05209_ VPWR VGND _05210_ sg13g2_a21oi_1
X_24937_ _04074_ _05202_ _05203_ _05210_ VPWR VGND 
+ _05211_
+ sg13g2_nor4_1
X_24938_ \atbs_core_0.spike_memory_0.n2417_o[15]\ _04623_ VPWR VGND _05212_ sg13g2_nor2_1
X_24939_ \atbs_core_0.spike_memory_0.n2414_o[15]\ _04702_ _03966_ VPWR VGND _05213_ sg13g2_o21ai_1
X_24940_ _04704_ _12590_ VPWR VGND _05214_ sg13g2_nor2_1
X_24941_ _12613_ _03852_ VPWR VGND _05215_ sg13g2_nor2_1
X_24942_ _04381_ _05214_ _05215_ _04343_ VPWR VGND 
+ _05216_
+ sg13g2_a22oi_1
X_24943_ _12590_ _04589_ VPWR VGND _05217_ sg13g2_nand2b_1
X_24944_ _04708_ _12613_ _05217_ VPWR VGND _05218_ sg13g2_o21ai_1
X_24945_ _03861_ _05218_ _03869_ VPWR VGND _05219_ sg13g2_a21oi_1
X_24946_ _04393_ _05216_ _05219_ VPWR VGND _05220_ sg13g2_a21oi_1
X_24947_ _05212_ _05213_ _05220_ VPWR VGND _05221_ sg13g2_nor3_1
X_24948_ \atbs_core_0.spike_memory_0.n2436_q[1212]\ _03804_ VPWR VGND _05222_ sg13g2_nor2_1
X_24949_ \atbs_core_0.spike_memory_0.n2418_o[15]\ _03946_ VPWR VGND _05223_ sg13g2_nor2_1
X_24950_ _03848_ _12648_ VPWR VGND _05224_ sg13g2_nor2_1
X_24951_ _12673_ _03852_ VPWR VGND _05225_ sg13g2_nor2_1
X_24952_ _04716_ _05224_ _05225_ _03857_ VPWR VGND 
+ _05226_
+ sg13g2_a22oi_1
X_24953_ _12648_ _03864_ VPWR VGND _05227_ sg13g2_nand2b_1
X_24954_ _04598_ _12673_ _05227_ VPWR VGND _05228_ sg13g2_o21ai_1
X_24955_ _03956_ _05228_ _04317_ VPWR VGND _05229_ sg13g2_a21oi_1
X_24956_ _03841_ _05226_ _05229_ VPWR VGND _05230_ sg13g2_a21oi_1
X_24957_ _12095_ _05222_ _05223_ _05230_ VPWR VGND 
+ _05231_
+ sg13g2_nor4_1
X_24958_ _05211_ _05221_ _05231_ VPWR VGND _05232_ sg13g2_nor3_1
X_24959_ \atbs_core_0.spike_memory_0.n2385_o[15]\ _03970_ VPWR VGND _05233_ sg13g2_nand2b_1
X_24960_ \atbs_core_0.spike_memory_0.n2382_o[15]\ _04771_ _05233_ VPWR VGND _05234_ sg13g2_o21ai_1
X_24961_ _03746_ _02305_ VPWR VGND _05235_ sg13g2_nor2_1
X_24962_ _02328_ _04006_ VPWR VGND _05236_ sg13g2_nor2_1
X_24963_ _03743_ _05235_ _05236_ _04512_ VPWR VGND 
+ _05237_
+ sg13g2_a22oi_1
X_24964_ _02305_ _04110_ VPWR VGND _05238_ sg13g2_nand2b_1
X_24965_ _04237_ _02328_ _05238_ VPWR VGND _05239_ sg13g2_o21ai_1
X_24966_ _04386_ _05239_ _04391_ VPWR VGND _05240_ sg13g2_a21oi_1
X_24967_ _04324_ _05237_ _05240_ VPWR VGND _05241_ sg13g2_a21oi_1
X_24968_ _05234_ _05241_ VPWR VGND _05242_ sg13g2_or2_1
X_24969_ \atbs_core_0.spike_memory_0.n2381_o[15]\ _12085_ VPWR VGND _05243_ sg13g2_nor2_1
X_24970_ \atbs_core_0.spike_memory_0.n2378_o[15]\ _04292_ VPWR VGND _05244_ sg13g2_nor2_1
X_24971_ _03741_ VPWR VGND _05245_ sg13g2_buf_1
X_24972_ _03854_ _02249_ VPWR VGND _05246_ sg13g2_nor2_1
X_24973_ _02273_ _03784_ VPWR VGND _05247_ sg13g2_nor2_1
X_24974_ _05245_ _05246_ _05247_ _03815_ VPWR VGND 
+ _05248_
+ sg13g2_a22oi_1
X_24975_ _02249_ _04455_ VPWR VGND _05249_ sg13g2_nand2b_1
X_24976_ _04050_ _02273_ _05249_ VPWR VGND _05250_ sg13g2_o21ai_1
X_24977_ _03757_ _05250_ _03867_ VPWR VGND _05251_ sg13g2_a21oi_1
X_24978_ _03992_ _05248_ _05251_ VPWR VGND _05252_ sg13g2_a21oi_1
X_24979_ _03773_ _05243_ _05244_ _05252_ VPWR VGND 
+ _05253_
+ sg13g2_nor4_1
X_24980_ \atbs_core_0.spike_memory_0.n2389_o[15]\ _03802_ VPWR VGND _05254_ sg13g2_nor2_1
X_24981_ \atbs_core_0.spike_memory_0.n2386_o[15]\ _04078_ VPWR VGND _05255_ sg13g2_nor2_1
X_24982_ _03988_ _02359_ VPWR VGND _05256_ sg13g2_nor2_1
X_24983_ _02382_ _03850_ VPWR VGND _05257_ sg13g2_nor2_1
X_24984_ _04062_ _05256_ _05257_ _04597_ VPWR VGND 
+ _05258_
+ sg13g2_a22oi_1
X_24985_ _02359_ _03981_ VPWR VGND _05259_ sg13g2_nand2b_1
X_24986_ _03846_ _02382_ _05259_ VPWR VGND _05260_ sg13g2_o21ai_1
X_24987_ _03859_ _05260_ _04068_ VPWR VGND _05261_ sg13g2_a21oi_1
X_24988_ _03839_ _05258_ _05261_ VPWR VGND _05262_ sg13g2_a21oi_1
X_24989_ _04746_ _05254_ _05255_ _05262_ VPWR VGND 
+ _05263_
+ sg13g2_nor4_1
X_24990_ _05253_ _05263_ _04276_ VPWR VGND _05264_ sg13g2_o21ai_1
X_24991_ _03924_ _05242_ _05264_ VPWR VGND _05265_ sg13g2_o21ai_1
X_24992_ \atbs_core_0.spike_memory_0.n2405_o[15]\ _04759_ VPWR VGND _05266_ sg13g2_nor2_1
X_24993_ \atbs_core_0.spike_memory_0.n2402_o[15]\ _03779_ VPWR VGND _05267_ sg13g2_nor2_1
X_24994_ _04254_ _02587_ VPWR VGND _05268_ sg13g2_nor2_1
X_24995_ _02608_ _03842_ VPWR VGND _05269_ sg13g2_nor2_1
X_24996_ _04108_ _05268_ _05269_ _03983_ VPWR VGND 
+ _05270_
+ sg13g2_a22oi_1
X_24997_ _02587_ _04088_ VPWR VGND _05271_ sg13g2_nand2b_1
X_24998_ _04425_ _02608_ _05271_ VPWR VGND _05272_ sg13g2_o21ai_1
X_24999_ _04010_ _05272_ _03810_ VPWR VGND _05273_ sg13g2_a21oi_1
X_25000_ _04118_ _05270_ _05273_ VPWR VGND _05274_ sg13g2_a21oi_1
X_25001_ _12093_ _05266_ _05267_ _05274_ VPWR VGND 
+ _05275_
+ sg13g2_nor4_1
X_25002_ \atbs_core_0.spike_memory_0.n2401_o[15]\ _12086_ VPWR VGND _05276_ sg13g2_nor2_1
X_25003_ \atbs_core_0.spike_memory_0.n2398_o[15]\ _04000_ _03780_ VPWR VGND _05277_ sg13g2_o21ai_1
X_25004_ _03787_ _02540_ VPWR VGND _05278_ sg13g2_nor2_1
X_25005_ _02561_ _03785_ VPWR VGND _05279_ sg13g2_nor2_1
X_25006_ _03782_ _05278_ _05279_ _03754_ VPWR VGND 
+ _05280_
+ sg13g2_a22oi_1
X_25007_ _02540_ _03891_ VPWR VGND _05281_ sg13g2_nand2b_1
X_25008_ _03753_ _02561_ _05281_ VPWR VGND _05282_ sg13g2_o21ai_1
X_25009_ _03758_ _05282_ _04294_ VPWR VGND _05283_ sg13g2_a21oi_1
X_25010_ _03739_ _05280_ _05283_ VPWR VGND _05284_ sg13g2_a21oi_1
X_25011_ _05276_ _05277_ _05284_ VPWR VGND _05285_ sg13g2_nor3_1
X_25012_ \atbs_core_0.spike_memory_0.n2397_o[15]\ _03876_ VPWR VGND _05286_ sg13g2_nor2_1
X_25013_ \atbs_core_0.spike_memory_0.n2394_o[15]\ _03835_ VPWR VGND _05287_ sg13g2_nor2_1
X_25014_ _04115_ _02492_ VPWR VGND _05288_ sg13g2_nor2_1
X_25015_ _02513_ _04006_ VPWR VGND _05289_ sg13g2_nor2_1
X_25016_ _04003_ _05288_ _05289_ _03978_ VPWR VGND 
+ _05290_
+ sg13g2_a22oi_1
X_25017_ _02492_ _04110_ VPWR VGND _05291_ sg13g2_nand2b_1
X_25018_ _03760_ _02513_ _05291_ VPWR VGND _05292_ sg13g2_o21ai_1
X_25019_ _04386_ _05292_ _04391_ VPWR VGND _05293_ sg13g2_a21oi_1
X_25020_ _04324_ _05290_ _05293_ VPWR VGND _05294_ sg13g2_a21oi_1
X_25021_ _03727_ _05286_ _05287_ _05294_ VPWR VGND 
+ _05295_
+ sg13g2_nor4_1
X_25022_ _05275_ _05285_ _05295_ VPWR VGND _05296_ sg13g2_or3_1
X_25023_ _03720_ _05265_ _05296_ _03717_ _04335_ VPWR 
+ VGND
+ _05297_ sg13g2_a221oi_1
X_25024_ _12079_ _05232_ _05297_ VPWR VGND _05298_ sg13g2_o21ai_1
X_25025_ _04503_ _05201_ _05298_ VPWR VGND _05299_ sg13g2_nand3_1
X_25026_ _04333_ _05174_ _05299_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[15]\ sg13g2_o21ai_1
X_25027_ \atbs_core_0.spike_memory_0.n2365_o[16]\ _04623_ VPWR VGND _05300_ sg13g2_nor2_1
X_25028_ \atbs_core_0.spike_memory_0.n2362_o[16]\ _04584_ VPWR VGND _05301_ sg13g2_nor2_1
X_25029_ _04590_ _12616_ VPWR VGND _05302_ sg13g2_nor2_1
X_25030_ _02017_ _03929_ VPWR VGND _05303_ sg13g2_nor2_1
X_25031_ _04588_ _05302_ _05303_ _04630_ VPWR VGND 
+ _05304_
+ sg13g2_a22oi_1
X_25032_ _12616_ _04598_ VPWR VGND _05305_ sg13g2_nand2b_1
X_25033_ _04593_ _02017_ _05305_ VPWR VGND _05306_ sg13g2_o21ai_1
X_25034_ _04596_ _05306_ _04635_ VPWR VGND _05307_ sg13g2_a21oi_1
X_25035_ _04626_ _05304_ _05307_ VPWR VGND _05308_ sg13g2_a21oi_1
X_25036_ _03872_ _05300_ _05301_ _05308_ VPWR VGND 
+ _05309_
+ sg13g2_nor4_1
X_25037_ \atbs_core_0.spike_memory_0.n2373_o[16]\ _04582_ VPWR VGND _05310_ sg13g2_nor2_1
X_25038_ \atbs_core_0.spike_memory_0.n2370_o[16]\ _04606_ VPWR VGND _05311_ sg13g2_nor2_1
X_25039_ _04610_ _02099_ VPWR VGND _05312_ sg13g2_nor2_1
X_25040_ _02122_ _03814_ VPWR VGND _05313_ sg13g2_nor2_1
X_25041_ _04609_ _05312_ _05313_ _04594_ VPWR VGND 
+ _05314_
+ sg13g2_a22oi_1
X_25042_ _02099_ _04708_ VPWR VGND _05315_ sg13g2_nand2b_1
X_25043_ _04616_ _02122_ _05315_ VPWR VGND _05316_ sg13g2_o21ai_1
X_25044_ _04615_ _05316_ _03812_ VPWR VGND _05317_ sg13g2_a21oi_1
X_25045_ _04586_ _05314_ _05317_ VPWR VGND _05318_ sg13g2_a21oi_1
X_25046_ _04219_ _05310_ _05311_ _05318_ VPWR VGND 
+ _05319_
+ sg13g2_nor4_1
X_25047_ _05309_ _05319_ _04504_ VPWR VGND _05320_ sg13g2_o21ai_1
X_25048_ \atbs_core_0.spike_memory_0.n2361_o[16]\ _04623_ VPWR VGND _05321_ sg13g2_nor2_1
X_25049_ \atbs_core_0.spike_memory_0.n2358_o[16]\ _03946_ VPWR VGND _05322_ sg13g2_nor2_1
X_25050_ _04593_ _02178_ VPWR VGND _05323_ sg13g2_nor2_1
X_25051_ _02340_ _04628_ VPWR VGND _05324_ sg13g2_nor2_1
X_25052_ _04662_ _05323_ _05324_ _04630_ VPWR VGND 
+ _05325_
+ sg13g2_a22oi_1
X_25053_ _02178_ _04052_ VPWR VGND _05326_ sg13g2_nand2b_1
X_25054_ _04632_ _02340_ _05326_ VPWR VGND _05327_ sg13g2_o21ai_1
X_25055_ _04666_ _05327_ _03880_ VPWR VGND _05328_ sg13g2_a21oi_1
X_25056_ _04626_ _05325_ _05328_ VPWR VGND _05329_ sg13g2_a21oi_1
X_25057_ _03872_ _05321_ _05322_ _05329_ VPWR VGND 
+ _05330_
+ sg13g2_nor4_1
X_25058_ \atbs_core_0.spike_memory_0.n2369_o[16]\ _04582_ VPWR VGND _05331_ sg13g2_nor2_1
X_25059_ \atbs_core_0.spike_memory_0.n2366_o[16]\ _04584_ VPWR VGND _05332_ sg13g2_nor2_1
X_25060_ _04616_ _02043_ VPWR VGND _05333_ sg13g2_nor2_1
X_25061_ _02065_ _03906_ VPWR VGND _05334_ sg13g2_nor2_1
X_25062_ _04588_ _05333_ _05334_ _04594_ VPWR VGND 
+ _05335_
+ sg13g2_a22oi_1
X_25063_ _02043_ _03856_ VPWR VGND _05336_ sg13g2_nand2b_1
X_25064_ _04590_ _02065_ _05336_ VPWR VGND _05337_ sg13g2_o21ai_1
X_25065_ _04596_ _05337_ _04149_ VPWR VGND _05338_ sg13g2_a21oi_1
X_25066_ _04586_ _05335_ _05338_ VPWR VGND _05339_ sg13g2_a21oi_1
X_25067_ _04219_ _05331_ _05332_ _05339_ VPWR VGND 
+ _05340_
+ sg13g2_nor4_1
X_25068_ _05330_ _05340_ _03725_ VPWR VGND _05341_ sg13g2_o21ai_1
X_25069_ _05320_ _05341_ VPWR VGND _05342_ sg13g2_and2_1
X_25070_ _04651_ _02408_ VPWR VGND _05343_ sg13g2_nor2_1
X_25071_ _02427_ _04510_ VPWR VGND _05344_ sg13g2_nor2_1
X_25072_ _04356_ _05343_ _05344_ _04680_ VPWR VGND 
+ _05345_
+ sg13g2_a22oi_1
X_25073_ _02408_ _04552_ VPWR VGND _05346_ sg13g2_nand2b_1
X_25074_ _04320_ _02427_ _05346_ VPWR VGND _05347_ sg13g2_o21ai_1
X_25075_ _04364_ _05347_ _04684_ VPWR VGND _05348_ sg13g2_a21oi_1
X_25076_ _04677_ _05345_ _05348_ VPWR VGND _05349_ sg13g2_a21oi_1
X_25077_ _00014_ _04675_ _04676_ _02466_ _05349_ VPWR 
+ VGND
+ _05350_ sg13g2_a221oi_1
X_25078_ _04632_ _02636_ VPWR VGND _05351_ sg13g2_nor2_1
X_25079_ _02657_ _03881_ VPWR VGND _05352_ sg13g2_nor2_1
X_25080_ _04662_ _05351_ _05352_ _04362_ VPWR VGND 
+ _05353_
+ sg13g2_a22oi_1
X_25081_ _02636_ _03957_ VPWR VGND _05354_ sg13g2_nand2b_1
X_25082_ _04365_ _02657_ _05354_ VPWR VGND _05355_ sg13g2_o21ai_1
X_25083_ _04666_ _05355_ _03880_ VPWR VGND _05356_ sg13g2_a21oi_1
X_25084_ _04355_ _05353_ _05356_ VPWR VGND _05357_ sg13g2_a21oi_1
X_25085_ _00013_ _04353_ _04354_ _02689_ _05357_ VPWR 
+ VGND
+ _05358_ sg13g2_a221oi_1
X_25086_ _04337_ _05350_ _05358_ _04673_ VPWR VGND 
+ _05359_
+ sg13g2_a22oi_1
X_25087_ _04651_ _02153_ VPWR VGND _05360_ sg13g2_nor2_1
X_25088_ _02176_ _03976_ VPWR VGND _05361_ sg13g2_nor2_1
X_25089_ _04339_ _05360_ _05361_ _04680_ VPWR VGND 
+ _05362_
+ sg13g2_a22oi_1
X_25090_ _02153_ _04552_ VPWR VGND _05363_ sg13g2_nand2b_1
X_25091_ _04340_ _02176_ _05363_ VPWR VGND _05364_ sg13g2_o21ai_1
X_25092_ _04345_ _05364_ _04684_ VPWR VGND _05365_ sg13g2_a21oi_1
X_25093_ _04677_ _05362_ _05365_ VPWR VGND _05366_ sg13g2_a21oi_1
X_25094_ _00015_ _04675_ _04676_ _02221_ _05366_ VPWR 
+ VGND
+ _05367_ sg13g2_a221oi_1
X_25095_ _04371_ _05367_ _04688_ VPWR VGND _05368_ sg13g2_a21oi_1
X_25096_ _05359_ _05368_ VPWR VGND _05369_ sg13g2_nand2_1
X_25097_ \atbs_core_0.spike_memory_0.n2413_o[16]\ _03901_ VPWR VGND _05370_ sg13g2_nor2_1
X_25098_ \atbs_core_0.spike_memory_0.n2410_o[16]\ _03903_ VPWR VGND _05371_ sg13g2_nor2_1
X_25099_ _03816_ _12536_ VPWR VGND _05372_ sg13g2_nor2_1
X_25100_ _12560_ _03819_ VPWR VGND _05373_ sg13g2_nor2_1
X_25101_ _04035_ _05372_ _05373_ _03911_ VPWR VGND 
+ _05374_
+ sg13g2_a22oi_1
X_25102_ _12536_ _03916_ VPWR VGND _05375_ sg13g2_nand2b_1
X_25103_ _03930_ _12560_ _05375_ VPWR VGND _05376_ sg13g2_o21ai_1
X_25104_ _03825_ _05376_ _04142_ VPWR VGND _05377_ sg13g2_a21oi_1
X_25105_ _03812_ _05374_ _05377_ VPWR VGND _05378_ sg13g2_a21oi_1
X_25106_ _04074_ _05370_ _05371_ _05378_ VPWR VGND 
+ _05379_
+ sg13g2_nor4_1
X_25107_ \atbs_core_0.spike_memory_0.n2417_o[16]\ _03804_ VPWR VGND _05380_ sg13g2_nor2_1
X_25108_ \atbs_core_0.spike_memory_0.n2414_o[16]\ _04702_ _03966_ VPWR VGND _05381_ sg13g2_o21ai_1
X_25109_ _04283_ _12591_ VPWR VGND _05382_ sg13g2_nor2_1
X_25110_ _12614_ _03852_ VPWR VGND _05383_ sg13g2_nor2_1
X_25111_ _04381_ _05382_ _05383_ _04343_ VPWR VGND 
+ _05384_
+ sg13g2_a22oi_1
X_25112_ _12591_ _04589_ VPWR VGND _05385_ sg13g2_nand2b_1
X_25113_ _04708_ _12614_ _05385_ VPWR VGND _05386_ sg13g2_o21ai_1
X_25114_ _03861_ _05386_ _03869_ VPWR VGND _05387_ sg13g2_a21oi_1
X_25115_ _04393_ _05384_ _05387_ VPWR VGND _05388_ sg13g2_a21oi_1
X_25116_ _05380_ _05381_ _05388_ VPWR VGND _05389_ sg13g2_nor3_1
X_25117_ \atbs_core_0.spike_memory_0.n2436_q[1213]\ _03804_ VPWR VGND _05390_ sg13g2_nor2_1
X_25118_ \atbs_core_0.spike_memory_0.n2418_o[16]\ _03946_ VPWR VGND _05391_ sg13g2_nor2_1
X_25119_ _03848_ _12649_ VPWR VGND _05392_ sg13g2_nor2_1
X_25120_ _12674_ _03852_ VPWR VGND _05393_ sg13g2_nor2_1
X_25121_ _04716_ _05392_ _05393_ _03857_ VPWR VGND 
+ _05394_
+ sg13g2_a22oi_1
X_25122_ _12649_ _03864_ VPWR VGND _05395_ sg13g2_nand2b_1
X_25123_ _04598_ _12674_ _05395_ VPWR VGND _05396_ sg13g2_o21ai_1
X_25124_ _03956_ _05396_ _04317_ VPWR VGND _05397_ sg13g2_a21oi_1
X_25125_ _03841_ _05394_ _05397_ VPWR VGND _05398_ sg13g2_a21oi_1
X_25126_ _12095_ _05390_ _05391_ _05398_ VPWR VGND 
+ _05399_
+ sg13g2_nor4_1
X_25127_ _05379_ _05389_ _05399_ VPWR VGND _05400_ sg13g2_nor3_1
X_25128_ \atbs_core_0.spike_memory_0.n2385_o[16]\ _03970_ VPWR VGND _05401_ sg13g2_nand2b_1
X_25129_ \atbs_core_0.spike_memory_0.n2382_o[16]\ _04771_ _05401_ VPWR VGND _05402_ sg13g2_o21ai_1
X_25130_ _03746_ _02306_ VPWR VGND _05403_ sg13g2_nor2_1
X_25131_ _02330_ _04006_ VPWR VGND _05404_ sg13g2_nor2_1
X_25132_ _03743_ _05403_ _05404_ _04512_ VPWR VGND 
+ _05405_
+ sg13g2_a22oi_1
X_25133_ _02306_ _04110_ VPWR VGND _05406_ sg13g2_nand2b_1
X_25134_ _04237_ _02330_ _05406_ VPWR VGND _05407_ sg13g2_o21ai_1
X_25135_ _04386_ _05407_ _04391_ VPWR VGND _05408_ sg13g2_a21oi_1
X_25136_ _04324_ _05405_ _05408_ VPWR VGND _05409_ sg13g2_a21oi_1
X_25137_ _05402_ _05409_ VPWR VGND _05410_ sg13g2_or2_1
X_25138_ \atbs_core_0.spike_memory_0.n2381_o[16]\ _12085_ VPWR VGND _05411_ sg13g2_nor2_1
X_25139_ \atbs_core_0.spike_memory_0.n2378_o[16]\ _04292_ VPWR VGND _05412_ sg13g2_nor2_1
X_25140_ _03854_ _02251_ VPWR VGND _05413_ sg13g2_nor2_1
X_25141_ _02274_ _03784_ VPWR VGND _05414_ sg13g2_nor2_1
X_25142_ _05245_ _05413_ _05414_ _03815_ VPWR VGND 
+ _05415_
+ sg13g2_a22oi_1
X_25143_ _02251_ _04455_ VPWR VGND _05416_ sg13g2_nand2b_1
X_25144_ _04050_ _02274_ _05416_ VPWR VGND _05417_ sg13g2_o21ai_1
X_25145_ _03757_ _05417_ _03867_ VPWR VGND _05418_ sg13g2_a21oi_1
X_25146_ _03992_ _05415_ _05418_ VPWR VGND _05419_ sg13g2_a21oi_1
X_25147_ _03726_ _05411_ _05412_ _05419_ VPWR VGND 
+ _05420_
+ sg13g2_nor4_1
X_25148_ \atbs_core_0.spike_memory_0.n2389_o[16]\ _03802_ VPWR VGND _05421_ sg13g2_nor2_1
X_25149_ \atbs_core_0.spike_memory_0.n2386_o[16]\ _04078_ VPWR VGND _05422_ sg13g2_nor2_1
X_25150_ _03988_ _02360_ VPWR VGND _05423_ sg13g2_nor2_1
X_25151_ _02383_ _03850_ VPWR VGND _05424_ sg13g2_nor2_1
X_25152_ _04062_ _05423_ _05424_ _04597_ VPWR VGND 
+ _05425_
+ sg13g2_a22oi_1
X_25153_ _02360_ _03981_ VPWR VGND _05426_ sg13g2_nand2b_1
X_25154_ _03846_ _02383_ _05426_ VPWR VGND _05427_ sg13g2_o21ai_1
X_25155_ _03859_ _05427_ _04068_ VPWR VGND _05428_ sg13g2_a21oi_1
X_25156_ _03839_ _05425_ _05428_ VPWR VGND _05429_ sg13g2_a21oi_1
X_25157_ _04746_ _05421_ _05422_ _05429_ VPWR VGND 
+ _05430_
+ sg13g2_nor4_1
X_25158_ _05420_ _05430_ _04276_ VPWR VGND _05431_ sg13g2_o21ai_1
X_25159_ _03924_ _05410_ _05431_ VPWR VGND _05432_ sg13g2_o21ai_1
X_25160_ \atbs_core_0.spike_memory_0.n2405_o[16]\ _04759_ VPWR VGND _05433_ sg13g2_nor2_1
X_25161_ \atbs_core_0.spike_memory_0.n2402_o[16]\ _03779_ VPWR VGND _05434_ sg13g2_nor2_1
X_25162_ _04254_ _02588_ VPWR VGND _05435_ sg13g2_nor2_1
X_25163_ _02609_ _03842_ VPWR VGND _05436_ sg13g2_nor2_1
X_25164_ _04108_ _05435_ _05436_ _03983_ VPWR VGND 
+ _05437_
+ sg13g2_a22oi_1
X_25165_ _02588_ _03988_ VPWR VGND _05438_ sg13g2_nand2b_1
X_25166_ _04425_ _02609_ _05438_ VPWR VGND _05439_ sg13g2_o21ai_1
X_25167_ _04010_ _05439_ _03810_ VPWR VGND _05440_ sg13g2_a21oi_1
X_25168_ _04118_ _05437_ _05440_ VPWR VGND _05441_ sg13g2_a21oi_1
X_25169_ _12093_ _05433_ _05434_ _05441_ VPWR VGND 
+ _05442_
+ sg13g2_nor4_1
X_25170_ \atbs_core_0.spike_memory_0.n2401_o[16]\ _12086_ VPWR VGND _05443_ sg13g2_nor2_1
X_25171_ \atbs_core_0.spike_memory_0.n2398_o[16]\ _04000_ _03722_ VPWR VGND _05444_ sg13g2_o21ai_1
X_25172_ _03787_ _02541_ VPWR VGND _05445_ sg13g2_nor2_1
X_25173_ _02562_ _03785_ VPWR VGND _05446_ sg13g2_nor2_1
X_25174_ _03782_ _05445_ _05446_ _03754_ VPWR VGND 
+ _05447_
+ sg13g2_a22oi_1
X_25175_ _02541_ _03891_ VPWR VGND _05448_ sg13g2_nand2b_1
X_25176_ _03753_ _02562_ _05448_ VPWR VGND _05449_ sg13g2_o21ai_1
X_25177_ _03758_ _05449_ _04294_ VPWR VGND _05450_ sg13g2_a21oi_1
X_25178_ _03739_ _05447_ _05450_ VPWR VGND _05451_ sg13g2_a21oi_1
X_25179_ _05443_ _05444_ _05451_ VPWR VGND _05452_ sg13g2_nor3_1
X_25180_ \atbs_core_0.spike_memory_0.n2397_o[16]\ _04759_ VPWR VGND _05453_ sg13g2_nor2_1
X_25181_ \atbs_core_0.spike_memory_0.n2394_o[16]\ _03835_ VPWR VGND _05454_ sg13g2_nor2_1
X_25182_ _04115_ _02493_ VPWR VGND _05455_ sg13g2_nor2_1
X_25183_ _02514_ _04006_ VPWR VGND _05456_ sg13g2_nor2_1
X_25184_ _04003_ _05455_ _05456_ _03978_ VPWR VGND 
+ _05457_
+ sg13g2_a22oi_1
X_25185_ _02493_ _04110_ VPWR VGND _05458_ sg13g2_nand2b_1
X_25186_ _04004_ _02514_ _05458_ VPWR VGND _05459_ sg13g2_o21ai_1
X_25187_ _04386_ _05459_ _04391_ VPWR VGND _05460_ sg13g2_a21oi_1
X_25188_ _04324_ _05457_ _05460_ VPWR VGND _05461_ sg13g2_a21oi_1
X_25189_ _03727_ _05453_ _05454_ _05461_ VPWR VGND 
+ _05462_
+ sg13g2_nor4_1
X_25190_ _05442_ _05452_ _05462_ VPWR VGND _05463_ sg13g2_or3_1
X_25191_ _03720_ _05432_ _05463_ _03717_ _04335_ VPWR 
+ VGND
+ _05464_ sg13g2_a221oi_1
X_25192_ _12079_ _05400_ _05464_ VPWR VGND _05465_ sg13g2_o21ai_1
X_25193_ _04503_ _05369_ _05465_ VPWR VGND _05466_ sg13g2_nand3_1
X_25194_ _04333_ _05342_ _05466_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[16]\ sg13g2_o21ai_1
X_25195_ _03984_ _02409_ VPWR VGND _05467_ sg13g2_nor2_1
X_25196_ _02428_ _03844_ VPWR VGND _05468_ sg13g2_nor2_1
X_25197_ _04609_ _05467_ _05468_ _04613_ VPWR VGND 
+ _05469_
+ sg13g2_a22oi_1
X_25198_ _02409_ _04704_ VPWR VGND _05470_ sg13g2_nand2b_1
X_25199_ _03984_ _02428_ _05470_ VPWR VGND _05471_ sg13g2_o21ai_1
X_25200_ _04615_ _05471_ _03948_ VPWR VGND _05472_ sg13g2_a21oi_1
X_25201_ _04608_ _05469_ _05472_ VPWR VGND _05473_ sg13g2_a21oi_1
X_25202_ _00017_ _04660_ _04661_ _02468_ _05473_ VPWR 
+ VGND
+ _05474_ sg13g2_a221oi_1
X_25203_ _04539_ _02637_ VPWR VGND _05475_ sg13g2_nor2_1
X_25204_ _02658_ _04555_ VPWR VGND _05476_ sg13g2_nor2_1
X_25205_ _04378_ _05475_ _05476_ _04384_ VPWR VGND 
+ _05477_
+ sg13g2_a22oi_1
X_25206_ _02637_ _04112_ VPWR VGND _05478_ sg13g2_nand2b_1
X_25207_ _04379_ _02658_ _05478_ VPWR VGND _05479_ sg13g2_o21ai_1
X_25208_ _04388_ _05479_ _04393_ VPWR VGND _05480_ sg13g2_a21oi_1
X_25209_ _04377_ _05477_ _05480_ VPWR VGND _05481_ sg13g2_a21oi_1
X_25210_ _00016_ _04660_ _04661_ _02691_ _05481_ VPWR 
+ VGND
+ _05482_ sg13g2_a221oi_1
X_25211_ _04673_ VPWR VGND _05483_ sg13g2_buf_1
X_25212_ _03718_ _05474_ _05482_ _05483_ VPWR VGND 
+ _05484_
+ sg13g2_a22oi_1
X_25213_ _03984_ _02155_ VPWR VGND _05485_ sg13g2_nor2_1
X_25214_ _02177_ _03844_ VPWR VGND _05486_ sg13g2_nor2_1
X_25215_ _04609_ _05485_ _05486_ _04613_ VPWR VGND 
+ _05487_
+ sg13g2_a22oi_1
X_25216_ _02155_ _04704_ VPWR VGND _05488_ sg13g2_nand2b_1
X_25217_ _04610_ _02177_ _05488_ VPWR VGND _05489_ sg13g2_o21ai_1
X_25218_ _04615_ _05489_ _03948_ VPWR VGND _05490_ sg13g2_a21oi_1
X_25219_ _04608_ _05487_ _05490_ VPWR VGND _05491_ sg13g2_a21oi_1
X_25220_ _00018_ _04660_ _04661_ _02223_ _05491_ VPWR 
+ VGND
+ _05492_ sg13g2_a221oi_1
X_25221_ _04330_ _05492_ _04688_ VPWR VGND _05493_ sg13g2_a21oi_1
X_25222_ \atbs_core_0.spike_memory_0.n2385_o[17]\ _03735_ VPWR VGND _05494_ sg13g2_nand2b_1
X_25223_ \atbs_core_0.spike_memory_0.n2382_o[17]\ _04102_ _05494_ VPWR VGND _05495_ sg13g2_o21ai_1
X_25224_ _03818_ VPWR VGND _05496_ sg13g2_buf_1
X_25225_ _04346_ _02307_ VPWR VGND _05497_ sg13g2_nor2_1
X_25226_ _02331_ _04265_ VPWR VGND _05498_ sg13g2_nor2_1
X_25227_ _05496_ _05497_ _05498_ _04112_ VPWR VGND 
+ _05499_
+ sg13g2_a22oi_1
X_25228_ _02307_ _03760_ VPWR VGND _05500_ sg13g2_nand2b_1
X_25229_ _04236_ _02331_ _05500_ VPWR VGND _05501_ sg13g2_o21ai_1
X_25230_ _04235_ _05501_ _03973_ VPWR VGND _05502_ sg13g2_a21oi_1
X_25231_ _03940_ _05499_ _05502_ VPWR VGND _05503_ sg13g2_a21oi_1
X_25232_ _05495_ _05503_ VPWR VGND _05504_ sg13g2_or2_1
X_25233_ \atbs_core_0.spike_memory_0.n2381_o[17]\ _04075_ VPWR VGND _05505_ sg13g2_nor2_1
X_25234_ \atbs_core_0.spike_memory_0.n2378_o[17]\ _04000_ VPWR VGND _05506_ sg13g2_nor2_1
X_25235_ _04480_ _02252_ VPWR VGND _05507_ sg13g2_nor2_1
X_25236_ _02275_ _05245_ VPWR VGND _05508_ sg13g2_nor2_1
X_25237_ _04422_ _05507_ _05508_ _04167_ VPWR VGND 
+ _05509_
+ sg13g2_a22oi_1
X_25238_ _04009_ VPWR VGND _05510_ sg13g2_buf_1
X_25239_ _02252_ _04050_ VPWR VGND _05511_ sg13g2_nand2b_1
X_25240_ _04054_ _02275_ _05511_ VPWR VGND _05512_ sg13g2_o21ai_1
X_25241_ _05510_ _05512_ _03738_ VPWR VGND _05513_ sg13g2_a21oi_1
X_25242_ _04839_ _05509_ _05513_ VPWR VGND _05514_ sg13g2_a21oi_1
X_25243_ _03773_ _05505_ _05506_ _05514_ VPWR VGND 
+ _05515_
+ sg13g2_nor4_1
X_25244_ \atbs_core_0.spike_memory_0.n2389_o[17]\ _04759_ VPWR VGND _05516_ sg13g2_nor2_1
X_25245_ \atbs_core_0.spike_memory_0.n2386_o[17]\ _04000_ VPWR VGND _05517_ sg13g2_nor2_1
X_25246_ _03863_ _02361_ VPWR VGND _05518_ sg13g2_nor2_1
X_25247_ _02385_ _05245_ VPWR VGND _05519_ sg13g2_nor2_1
X_25248_ _04250_ _05518_ _05519_ _03864_ VPWR VGND 
+ _05520_
+ sg13g2_a22oi_1
X_25249_ _02361_ _03846_ VPWR VGND _05521_ sg13g2_nand2b_1
X_25250_ _03863_ _02385_ _05521_ VPWR VGND _05522_ sg13g2_o21ai_1
X_25251_ _05510_ _05522_ _03810_ VPWR VGND _05523_ sg13g2_a21oi_1
X_25252_ _04098_ _05520_ _05523_ VPWR VGND _05524_ sg13g2_a21oi_1
X_25253_ _04746_ _05516_ _05517_ _05524_ VPWR VGND 
+ _05525_
+ sg13g2_nor4_1
X_25254_ _05515_ _05525_ _03924_ VPWR VGND _05526_ sg13g2_o21ai_1
X_25255_ _04277_ _05504_ _05526_ VPWR VGND _05527_ sg13g2_o21ai_1
X_25256_ \atbs_core_0.spike_memory_0.n2405_o[17]\ _04245_ VPWR VGND _05528_ sg13g2_nor2_1
X_25257_ \atbs_core_0.spike_memory_0.n2402_o[17]\ _04247_ VPWR VGND _05529_ sg13g2_nor2_1
X_25258_ _04413_ _02589_ VPWR VGND _05530_ sg13g2_nor2_1
X_25259_ _02610_ _04086_ VPWR VGND _05531_ sg13g2_nor2_1
X_25260_ _03751_ _05530_ _05531_ _04704_ VPWR VGND 
+ _05532_
+ sg13g2_a22oi_1
X_25261_ _03988_ VPWR VGND _05533_ sg13g2_buf_1
X_25262_ _02589_ _04425_ VPWR VGND _05534_ sg13g2_nand2b_1
X_25263_ _05533_ _02610_ _05534_ VPWR VGND _05535_ sg13g2_o21ai_1
X_25264_ _04092_ _05535_ _04839_ VPWR VGND _05536_ sg13g2_a21oi_1
X_25265_ _03769_ _05532_ _05536_ VPWR VGND _05537_ sg13g2_a21oi_1
X_25266_ _12094_ _05528_ _05529_ _05537_ VPWR VGND 
+ _05538_
+ sg13g2_nor4_1
X_25267_ \atbs_core_0.spike_memory_0.n2401_o[17]\ _04372_ VPWR VGND _05539_ sg13g2_nor2_1
X_25268_ _04292_ VPWR VGND _05540_ sg13g2_buf_1
X_25269_ \atbs_core_0.spike_memory_0.n2398_o[17]\ _05540_ _03723_ VPWR VGND _05541_ sg13g2_o21ai_1
X_25270_ _04026_ _02542_ VPWR VGND _05542_ sg13g2_nor2_1
X_25271_ _02563_ _03975_ VPWR VGND _05543_ sg13g2_nor2_1
X_25272_ _04105_ VPWR VGND _05544_ sg13g2_buf_1
X_25273_ _04152_ _05542_ _05543_ _05544_ VPWR VGND 
+ _05545_
+ sg13g2_a22oi_1
X_25274_ _02542_ _03753_ VPWR VGND _05546_ sg13g2_nand2b_1
X_25275_ _03764_ _02563_ _05546_ VPWR VGND _05547_ sg13g2_o21ai_1
X_25276_ _04114_ _05547_ _04118_ VPWR VGND _05548_ sg13g2_a21oi_1
X_25277_ _04142_ _05545_ _05548_ VPWR VGND _05549_ sg13g2_a21oi_1
X_25278_ _05539_ _05541_ _05549_ VPWR VGND _05550_ sg13g2_nor3_1
X_25279_ \atbs_core_0.spike_memory_0.n2397_o[17]\ _04260_ VPWR VGND _05551_ sg13g2_nor2_1
X_25280_ \atbs_core_0.spike_memory_0.n2394_o[17]\ _04079_ VPWR VGND _05552_ sg13g2_nor2_1
X_25281_ _04111_ _02495_ VPWR VGND _05553_ sg13g2_nor2_1
X_25282_ _02516_ _04265_ VPWR VGND _05554_ sg13g2_nor2_1
X_25283_ _03884_ _05553_ _05554_ _04268_ VPWR VGND 
+ _05555_
+ sg13g2_a22oi_1
X_25284_ _02495_ _04004_ VPWR VGND _05556_ sg13g2_nand2b_1
X_25285_ _04083_ _02516_ _05556_ VPWR VGND _05557_ sg13g2_o21ai_1
X_25286_ _04253_ _05557_ _04272_ VPWR VGND _05558_ sg13g2_a21oi_1
X_25287_ _04263_ _05555_ _05558_ VPWR VGND _05559_ sg13g2_a21oi_1
X_25288_ _03774_ _05551_ _05552_ _05559_ VPWR VGND 
+ _05560_
+ sg13g2_nor4_1
X_25289_ _05538_ _05550_ _05560_ VPWR VGND _05561_ sg13g2_or3_1
X_25290_ _04330_ _05527_ _05561_ _03718_ _04336_ VPWR 
+ VGND
+ _05562_ sg13g2_a221oi_1
X_25291_ \atbs_core_0.spike_memory_0.n2413_o[17]\ _03803_ VPWR VGND _05563_ sg13g2_nor2_1
X_25292_ \atbs_core_0.spike_memory_0.n2410_o[17]\ _05540_ VPWR VGND _05564_ sg13g2_nor2_1
X_25293_ _04597_ _12538_ VPWR VGND _05565_ sg13g2_nor2_1
X_25294_ _12561_ _03851_ VPWR VGND _05566_ sg13g2_nor2_1
X_25295_ _03843_ _05565_ _05566_ _03949_ VPWR VGND 
+ _05567_
+ sg13g2_a22oi_1
X_25296_ _12538_ _04480_ VPWR VGND _05568_ sg13g2_nand2b_1
X_25297_ _04051_ _12561_ _05568_ VPWR VGND _05569_ sg13g2_o21ai_1
X_25298_ _03955_ _05569_ _03868_ VPWR VGND _05570_ sg13g2_a21oi_1
X_25299_ _03993_ _05567_ _05570_ VPWR VGND _05571_ sg13g2_a21oi_1
X_25300_ _04244_ _05563_ _05564_ _05571_ VPWR VGND 
+ _05572_
+ sg13g2_nor4_1
X_25301_ \atbs_core_0.spike_memory_0.n2436_q[1214]\ _03803_ VPWR VGND _05573_ sg13g2_nor2_1
X_25302_ \atbs_core_0.spike_memory_0.n2418_o[17]\ _05540_ VPWR VGND _05574_ sg13g2_nor2_1
X_25303_ _03847_ _12650_ VPWR VGND _05575_ sg13g2_nor2_1
X_25304_ _12675_ _03851_ VPWR VGND _05576_ sg13g2_nor2_1
X_25305_ _03843_ _05575_ _05576_ _03848_ VPWR VGND 
+ _05577_
+ sg13g2_a22oi_1
X_25306_ _12650_ _03982_ VPWR VGND _05578_ sg13g2_nand2b_1
X_25307_ _04597_ _12675_ _05578_ VPWR VGND _05579_ sg13g2_o21ai_1
X_25308_ _03860_ _05579_ _04287_ VPWR VGND _05580_ sg13g2_a21oi_1
X_25309_ _03840_ _05577_ _05580_ VPWR VGND _05581_ sg13g2_a21oi_1
X_25310_ _03899_ _05573_ _05574_ _05581_ VPWR VGND 
+ _05582_
+ sg13g2_nor4_1
X_25311_ _05572_ _05582_ _04277_ VPWR VGND _05583_ sg13g2_o21ai_1
X_25312_ _05583_ VPWR VGND _05584_ sg13g2_inv_1
X_25313_ \atbs_core_0.spike_memory_0.n2417_o[17]\ _03736_ VPWR VGND _05585_ sg13g2_nand2b_1
X_25314_ \atbs_core_0.spike_memory_0.n2414_o[17]\ _03946_ _05585_ VPWR VGND _05586_ sg13g2_o21ai_1
X_25315_ _04383_ _12593_ VPWR VGND _05587_ sg13g2_nor2_1
X_25316_ _12615_ _03844_ VPWR VGND _05588_ sg13g2_nor2_1
X_25317_ _04609_ _05587_ _05588_ _04613_ VPWR VGND 
+ _05589_
+ sg13g2_a22oi_1
X_25318_ _12593_ _04090_ VPWR VGND _05590_ sg13g2_nand2b_1
X_25319_ _03984_ _12615_ _05590_ VPWR VGND _05591_ sg13g2_o21ai_1
X_25320_ _04615_ _05591_ _03841_ VPWR VGND _05592_ sg13g2_a21oi_1
X_25321_ _04608_ _05589_ _05592_ VPWR VGND _05593_ sg13g2_a21oi_1
X_25322_ _03925_ _04604_ _05586_ _05593_ VPWR VGND 
+ _05594_
+ sg13g2_nor4_1
X_25323_ _05584_ _05594_ _05483_ VPWR VGND _05595_ sg13g2_o21ai_1
X_25324_ _05484_ _05493_ _05562_ _05595_ VPWR VGND 
+ _05596_
+ sg13g2_a22oi_1
X_25325_ \atbs_core_0.spike_memory_0.n2361_o[17]\ _04506_ VPWR VGND _05597_ sg13g2_nor2_1
X_25326_ \atbs_core_0.spike_memory_0.n2358_o[17]\ _04508_ VPWR VGND _05598_ sg13g2_nor2_1
X_25327_ _04513_ _02202_ VPWR VGND _05599_ sg13g2_nor2_1
X_25328_ _02352_ _04716_ VPWR VGND _05600_ sg13g2_nor2_1
X_25329_ _04511_ _05599_ _05600_ _04384_ VPWR VGND 
+ _05601_
+ sg13g2_a22oi_1
X_25330_ _02202_ _04518_ VPWR VGND _05602_ sg13g2_nand2b_1
X_25331_ _04383_ _02352_ _05602_ VPWR VGND _05603_ sg13g2_o21ai_1
X_25332_ _04517_ _05603_ _04521_ VPWR VGND _05604_ sg13g2_a21oi_1
X_25333_ _04377_ _05601_ _05604_ VPWR VGND _05605_ sg13g2_a21oi_1
X_25334_ _04505_ _05597_ _05598_ _05605_ VPWR VGND 
+ _05606_
+ sg13g2_nor4_1
X_25335_ \atbs_core_0.spike_memory_0.n2369_o[17]\ _04525_ VPWR VGND _05607_ sg13g2_nor2_1
X_25336_ \atbs_core_0.spike_memory_0.n2366_o[17]\ _04549_ VPWR VGND _05608_ sg13g2_nor2_1
X_25337_ _04553_ _02044_ VPWR VGND _05609_ sg13g2_nor2_1
X_25338_ _02066_ _04533_ VPWR VGND _05610_ sg13g2_nor2_1
X_25339_ _04531_ _05609_ _05610_ _04536_ VPWR VGND 
+ _05611_
+ sg13g2_a22oi_1
X_25340_ _02044_ _04559_ VPWR VGND _05612_ sg13g2_nand2b_1
X_25341_ _04539_ _02066_ _05612_ VPWR VGND _05613_ sg13g2_o21ai_1
X_25342_ _04538_ _05613_ _04542_ VPWR VGND _05614_ sg13g2_a21oi_1
X_25343_ _04530_ _05611_ _05614_ VPWR VGND _05615_ sg13g2_a21oi_1
X_25344_ _04604_ _05607_ _05608_ _05615_ VPWR VGND 
+ _05616_
+ sg13g2_nor4_1
X_25345_ _04504_ _05606_ _05616_ VPWR VGND _05617_ sg13g2_nor3_1
X_25346_ \atbs_core_0.spike_memory_0.n2365_o[17]\ _04506_ VPWR VGND _05618_ sg13g2_nor2_1
X_25347_ \atbs_core_0.spike_memory_0.n2362_o[17]\ _04549_ VPWR VGND _05619_ sg13g2_nor2_1
X_25348_ _04553_ _12619_ VPWR VGND _05620_ sg13g2_nor2_1
X_25349_ _02018_ _04555_ VPWR VGND _05621_ sg13g2_nor2_1
X_25350_ _04378_ _05620_ _05621_ _04557_ VPWR VGND 
+ _05622_
+ sg13g2_a22oi_1
X_25351_ _12619_ _04559_ VPWR VGND _05623_ sg13g2_nand2b_1
X_25352_ _03755_ _02018_ _05623_ VPWR VGND _05624_ sg13g2_o21ai_1
X_25353_ _04388_ _05624_ _04562_ VPWR VGND _05625_ sg13g2_a21oi_1
X_25354_ _04551_ _05622_ _05625_ VPWR VGND _05626_ sg13g2_a21oi_1
X_25355_ _03729_ _05618_ _05619_ _05626_ VPWR VGND 
+ _05627_
+ sg13g2_nor4_1
X_25356_ \atbs_core_0.spike_memory_0.n2373_o[17]\ _12088_ VPWR VGND _05628_ sg13g2_nor2_1
X_25357_ \atbs_core_0.spike_memory_0.n2370_o[17]\ _04528_ VPWR VGND _05629_ sg13g2_nor2_1
X_25358_ _03934_ _02100_ VPWR VGND _05630_ sg13g2_nor2_1
X_25359_ _02123_ _04570_ VPWR VGND _05631_ sg13g2_nor2_1
X_25360_ _04568_ _05630_ _05631_ _02714_ VPWR VGND 
+ _05632_
+ sg13g2_a22oi_1
X_25361_ _02100_ _04361_ VPWR VGND _05633_ sg13g2_nand2b_1
X_25362_ _04574_ _02123_ _05633_ VPWR VGND _05634_ sg13g2_o21ai_1
X_25363_ _04573_ _05634_ _04338_ VPWR VGND _05635_ sg13g2_a21oi_1
X_25364_ _02702_ _05632_ _05635_ VPWR VGND _05636_ sg13g2_a21oi_1
X_25365_ _04126_ _05628_ _05629_ _05636_ VPWR VGND 
+ _05637_
+ sg13g2_nor4_1
X_25366_ _04547_ _05627_ _05637_ VPWR VGND _05638_ sg13g2_nor3_1
X_25367_ _07549_ _05617_ _05638_ VPWR VGND _05639_ sg13g2_nor3_1
X_25368_ _04333_ _05596_ _05639_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[17]\ sg13g2_a21o_1
X_25369_ _04340_ _02410_ VPWR VGND _05640_ sg13g2_nor2_1
X_25370_ _02429_ _03976_ VPWR VGND _05641_ sg13g2_nor2_1
X_25371_ _04339_ _05640_ _05641_ _04680_ VPWR VGND 
+ _05642_
+ sg13g2_a22oi_1
X_25372_ _02410_ _03788_ VPWR VGND _05643_ sg13g2_nand2b_1
X_25373_ _04347_ _02429_ _05643_ VPWR VGND _05644_ sg13g2_o21ai_1
X_25374_ _04345_ _05644_ _04684_ VPWR VGND _05645_ sg13g2_a21oi_1
X_25375_ _04677_ _05642_ _05645_ VPWR VGND _05646_ sg13g2_a21oi_1
X_25376_ _00020_ _04675_ _04676_ _02470_ _05646_ VPWR 
+ VGND
+ _05647_ sg13g2_a221oi_1
X_25377_ _04357_ _02156_ VPWR VGND _05648_ sg13g2_nor2_1
X_25378_ _02179_ _03881_ VPWR VGND _05649_ sg13g2_nor2_1
X_25379_ _04662_ _05648_ _05649_ _04362_ VPWR VGND 
+ _05650_
+ sg13g2_a22oi_1
X_25380_ _02156_ _03816_ VPWR VGND _05651_ sg13g2_nand2b_1
X_25381_ _04365_ _02179_ _05651_ VPWR VGND _05652_ sg13g2_o21ai_1
X_25382_ _04666_ _05652_ _04021_ VPWR VGND _05653_ sg13g2_a21oi_1
X_25383_ _04355_ _05650_ _05653_ VPWR VGND _05654_ sg13g2_a21oi_1
X_25384_ _00021_ _04353_ _04354_ _02225_ _05654_ VPWR 
+ VGND
+ _05655_ sg13g2_a221oi_1
X_25385_ _04337_ _05647_ _05655_ _04330_ _04688_ VPWR 
+ VGND
+ _05656_ sg13g2_a221oi_1
X_25386_ _02713_ _02638_ VPWR VGND _05657_ sg13g2_nor2_1
X_25387_ _02659_ _04570_ VPWR VGND _05658_ sg13g2_nor2_1
X_25388_ _04568_ _05657_ _05658_ _04536_ VPWR VGND 
+ _05659_
+ sg13g2_a22oi_1
X_25389_ _02638_ _04320_ VPWR VGND _05660_ sg13g2_nand2b_1
X_25390_ _04574_ _02659_ _05660_ VPWR VGND _05661_ sg13g2_o21ai_1
X_25391_ _04573_ _05661_ _04542_ VPWR VGND _05662_ sg13g2_a21oi_1
X_25392_ _04530_ _05659_ _05662_ VPWR VGND _05663_ sg13g2_a21oi_1
X_25393_ _00019_ _04660_ _04661_ _02693_ _05663_ VPWR 
+ VGND
+ _05664_ sg13g2_a221oi_1
X_25394_ _05483_ _05664_ VPWR VGND _05665_ sg13g2_nand2_1
X_25395_ \atbs_core_0.spike_memory_0.n2385_o[18]\ _03735_ VPWR VGND _05666_ sg13g2_nand2b_1
X_25396_ \atbs_core_0.spike_memory_0.n2382_o[18]\ _04102_ _05666_ VPWR VGND _05667_ sg13g2_o21ai_1
X_25397_ _04346_ _02308_ VPWR VGND _05668_ sg13g2_nor2_1
X_25398_ _02332_ _04265_ VPWR VGND _05669_ sg13g2_nor2_1
X_25399_ _05496_ _05668_ _05669_ _04112_ VPWR VGND 
+ _05670_
+ sg13g2_a22oi_1
X_25400_ _02308_ _03760_ VPWR VGND _05671_ sg13g2_nand2b_1
X_25401_ _04236_ _02332_ _05671_ VPWR VGND _05672_ sg13g2_o21ai_1
X_25402_ _04235_ _05672_ _03973_ VPWR VGND _05673_ sg13g2_a21oi_1
X_25403_ _03940_ _05670_ _05673_ VPWR VGND _05674_ sg13g2_a21oi_1
X_25404_ _05667_ _05674_ VPWR VGND _05675_ sg13g2_or2_1
X_25405_ \atbs_core_0.spike_memory_0.n2381_o[18]\ _04075_ VPWR VGND _05676_ sg13g2_nor2_1
X_25406_ \atbs_core_0.spike_memory_0.n2378_o[18]\ _04229_ VPWR VGND _05677_ sg13g2_nor2_1
X_25407_ _04480_ _02253_ VPWR VGND _05678_ sg13g2_nor2_1
X_25408_ _02276_ _03742_ VPWR VGND _05679_ sg13g2_nor2_1
X_25409_ _04422_ _05678_ _05679_ _03827_ VPWR VGND 
+ _05680_
+ sg13g2_a22oi_1
X_25410_ _02253_ _04050_ VPWR VGND _05681_ sg13g2_nand2b_1
X_25411_ _03915_ _02276_ _05681_ VPWR VGND _05682_ sg13g2_o21ai_1
X_25412_ _05510_ _05682_ _03738_ VPWR VGND _05683_ sg13g2_a21oi_1
X_25413_ _04839_ _05680_ _05683_ VPWR VGND _05684_ sg13g2_a21oi_1
X_25414_ _03773_ _05676_ _05677_ _05684_ VPWR VGND 
+ _05685_
+ sg13g2_nor4_1
X_25415_ \atbs_core_0.spike_memory_0.n2389_o[18]\ _04759_ VPWR VGND _05686_ sg13g2_nor2_1
X_25416_ \atbs_core_0.spike_memory_0.n2386_o[18]\ _04000_ VPWR VGND _05687_ sg13g2_nor2_1
X_25417_ _03863_ _02364_ VPWR VGND _05688_ sg13g2_nor2_1
X_25418_ _02386_ _05245_ VPWR VGND _05689_ sg13g2_nor2_1
X_25419_ _04250_ _05688_ _05689_ _03864_ VPWR VGND 
+ _05690_
+ sg13g2_a22oi_1
X_25420_ _02364_ _03846_ VPWR VGND _05691_ sg13g2_nand2b_1
X_25421_ _03863_ _02386_ _05691_ VPWR VGND _05692_ sg13g2_o21ai_1
X_25422_ _05510_ _05692_ _03810_ VPWR VGND _05693_ sg13g2_a21oi_1
X_25423_ _04098_ _05690_ _05693_ VPWR VGND _05694_ sg13g2_a21oi_1
X_25424_ _04746_ _05686_ _05687_ _05694_ VPWR VGND 
+ _05695_
+ sg13g2_nor4_1
X_25425_ _05685_ _05695_ _03924_ VPWR VGND _05696_ sg13g2_o21ai_1
X_25426_ _04277_ _05675_ _05696_ VPWR VGND _05697_ sg13g2_o21ai_1
X_25427_ \atbs_core_0.spike_memory_0.n2405_o[18]\ _04245_ VPWR VGND _05698_ sg13g2_nor2_1
X_25428_ \atbs_core_0.spike_memory_0.n2402_o[18]\ _04247_ VPWR VGND _05699_ sg13g2_nor2_1
X_25429_ _04413_ _02590_ VPWR VGND _05700_ sg13g2_nor2_1
X_25430_ _02612_ _04086_ VPWR VGND _05701_ sg13g2_nor2_1
X_25431_ _04280_ _05700_ _05701_ _04704_ VPWR VGND 
+ _05702_
+ sg13g2_a22oi_1
X_25432_ _02590_ _04425_ VPWR VGND _05703_ sg13g2_nand2b_1
X_25433_ _05533_ _02612_ _05703_ VPWR VGND _05704_ sg13g2_o21ai_1
X_25434_ _04092_ _05704_ _04839_ VPWR VGND _05705_ sg13g2_a21oi_1
X_25435_ _03769_ _05702_ _05705_ VPWR VGND _05706_ sg13g2_a21oi_1
X_25436_ _12094_ _05698_ _05699_ _05706_ VPWR VGND 
+ _05707_
+ sg13g2_nor4_1
X_25437_ \atbs_core_0.spike_memory_0.n2401_o[18]\ _04372_ VPWR VGND _05708_ sg13g2_nor2_1
X_25438_ \atbs_core_0.spike_memory_0.n2398_o[18]\ _05540_ _03723_ VPWR VGND _05709_ sg13g2_o21ai_1
X_25439_ _04026_ _02543_ VPWR VGND _05710_ sg13g2_nor2_1
X_25440_ _02564_ _03975_ VPWR VGND _05711_ sg13g2_nor2_1
X_25441_ _04152_ _05710_ _05711_ _05544_ VPWR VGND 
+ _05712_
+ sg13g2_a22oi_1
X_25442_ _02543_ _04115_ VPWR VGND _05713_ sg13g2_nand2b_1
X_25443_ _03764_ _02564_ _05713_ VPWR VGND _05714_ sg13g2_o21ai_1
X_25444_ _04114_ _05714_ _04118_ VPWR VGND _05715_ sg13g2_a21oi_1
X_25445_ _04142_ _05712_ _05715_ VPWR VGND _05716_ sg13g2_a21oi_1
X_25446_ _05708_ _05709_ _05716_ VPWR VGND _05717_ sg13g2_nor3_1
X_25447_ \atbs_core_0.spike_memory_0.n2397_o[18]\ _04260_ VPWR VGND _05718_ sg13g2_nor2_1
X_25448_ \atbs_core_0.spike_memory_0.n2394_o[18]\ _04079_ VPWR VGND _05719_ sg13g2_nor2_1
X_25449_ _04236_ _02496_ VPWR VGND _05720_ sg13g2_nor2_1
X_25450_ _02517_ _04265_ VPWR VGND _05721_ sg13g2_nor2_1
X_25451_ _03884_ _05720_ _05721_ _04268_ VPWR VGND 
+ _05722_
+ sg13g2_a22oi_1
X_25452_ _02496_ _04004_ VPWR VGND _05723_ sg13g2_nand2b_1
X_25453_ _04083_ _02517_ _05723_ VPWR VGND _05724_ sg13g2_o21ai_1
X_25454_ _04253_ _05724_ _04272_ VPWR VGND _05725_ sg13g2_a21oi_1
X_25455_ _04263_ _05722_ _05725_ VPWR VGND _05726_ sg13g2_a21oi_1
X_25456_ _04244_ _05718_ _05719_ _05726_ VPWR VGND 
+ _05727_
+ sg13g2_nor4_1
X_25457_ _05707_ _05717_ _05727_ VPWR VGND _05728_ sg13g2_or3_1
X_25458_ _04330_ _05697_ _05728_ _03718_ _04336_ VPWR 
+ VGND
+ _05729_ sg13g2_a221oi_1
X_25459_ \atbs_core_0.spike_memory_0.n2413_o[18]\ _04372_ VPWR VGND _05730_ sg13g2_nor2_1
X_25460_ \atbs_core_0.spike_memory_0.n2410_o[18]\ _04527_ VPWR VGND _05731_ sg13g2_nor2_1
X_25461_ _03747_ _12539_ VPWR VGND _05732_ sg13g2_nor2_1
X_25462_ _12562_ _03751_ VPWR VGND _05733_ sg13g2_nor2_1
X_25463_ _03744_ _05732_ _05733_ _04379_ VPWR VGND 
+ _05734_
+ sg13g2_a22oi_1
X_25464_ _12539_ _03764_ VPWR VGND _05735_ sg13g2_nand2b_1
X_25465_ _04512_ _12562_ _05735_ VPWR VGND _05736_ sg13g2_o21ai_1
X_25466_ _03759_ _05736_ _04392_ VPWR VGND _05737_ sg13g2_a21oi_1
X_25467_ _03740_ _05734_ _05737_ VPWR VGND _05738_ sg13g2_a21oi_1
X_25468_ _03800_ _05730_ _05731_ _05738_ VPWR VGND 
+ _05739_
+ sg13g2_nor4_1
X_25469_ \atbs_core_0.spike_memory_0.n2417_o[18]\ _03944_ VPWR VGND _05740_ sg13g2_nor2_1
X_25470_ \atbs_core_0.spike_memory_0.n2414_o[18]\ _04032_ _03966_ VPWR VGND _05741_ sg13g2_o21ai_1
X_25471_ _03907_ _12594_ VPWR VGND _05742_ sg13g2_nor2_1
X_25472_ _12617_ _03909_ VPWR VGND _05743_ sg13g2_nor2_1
X_25473_ _03906_ _05742_ _05743_ _03911_ VPWR VGND 
+ _05744_
+ sg13g2_a22oi_1
X_25474_ _03791_ VPWR VGND _05745_ sg13g2_buf_1
X_25475_ _12594_ _05745_ VPWR VGND _05746_ sg13g2_nand2b_1
X_25476_ _03914_ _12617_ _05746_ VPWR VGND _05747_ sg13g2_o21ai_1
X_25477_ _03913_ _05747_ _03919_ VPWR VGND _05748_ sg13g2_a21oi_1
X_25478_ _03905_ _05744_ _05748_ VPWR VGND _05749_ sg13g2_a21oi_1
X_25479_ _05740_ _05741_ _05749_ VPWR VGND _05750_ sg13g2_nor3_1
X_25480_ \atbs_core_0.spike_memory_0.n2436_q[1215]\ _03877_ VPWR VGND _05751_ sg13g2_nor2_1
X_25481_ \atbs_core_0.spike_memory_0.n2418_o[18]\ _04702_ VPWR VGND _05752_ sg13g2_nor2_1
X_25482_ _03821_ VPWR VGND _05753_ sg13g2_buf_1
X_25483_ _05753_ _12651_ VPWR VGND _05754_ sg13g2_nor2_1
X_25484_ _12677_ _05496_ VPWR VGND _05755_ sg13g2_nor2_1
X_25485_ _03929_ _05754_ _05755_ _02713_ VPWR VGND 
+ _05756_
+ sg13g2_a22oi_1
X_25486_ _12651_ _03892_ VPWR VGND _05757_ sg13g2_nand2b_1
X_25487_ _02712_ _12677_ _05757_ VPWR VGND _05758_ sg13g2_o21ai_1
X_25488_ _03889_ _05758_ _04263_ VPWR VGND _05759_ sg13g2_a21oi_1
X_25489_ _04635_ _05756_ _05759_ VPWR VGND _05760_ sg13g2_a21oi_1
X_25490_ _12095_ _05751_ _05752_ _05760_ VPWR VGND 
+ _05761_
+ sg13g2_nor4_1
X_25491_ _05739_ _05750_ _05761_ VPWR VGND _05762_ sg13g2_nor3_1
X_25492_ _05762_ _05483_ VPWR VGND _05763_ sg13g2_nand2b_1
X_25493_ _05656_ _05665_ _05729_ _05763_ VPWR VGND 
+ _05764_
+ sg13g2_a22oi_1
X_25494_ \atbs_core_0.spike_memory_0.n2361_o[18]\ _04506_ VPWR VGND _05765_ sg13g2_nor2_1
X_25495_ \atbs_core_0.spike_memory_0.n2358_o[18]\ _04508_ VPWR VGND _05766_ sg13g2_nor2_1
X_25496_ _04513_ _02227_ VPWR VGND _05767_ sg13g2_nor2_1
X_25497_ _02365_ _04716_ VPWR VGND _05768_ sg13g2_nor2_1
X_25498_ _04511_ _05767_ _05768_ _04384_ VPWR VGND 
+ _05769_
+ sg13g2_a22oi_1
X_25499_ _02227_ _04518_ VPWR VGND _05770_ sg13g2_nand2b_1
X_25500_ _04383_ _02365_ _05770_ VPWR VGND _05771_ sg13g2_o21ai_1
X_25501_ _04517_ _05771_ _04521_ VPWR VGND _05772_ sg13g2_a21oi_1
X_25502_ _04377_ _05769_ _05772_ VPWR VGND _05773_ sg13g2_a21oi_1
X_25503_ _04505_ _05765_ _05766_ _05773_ VPWR VGND 
+ _05774_
+ sg13g2_nor4_1
X_25504_ \atbs_core_0.spike_memory_0.n2369_o[18]\ _04525_ VPWR VGND _05775_ sg13g2_nor2_1
X_25505_ \atbs_core_0.spike_memory_0.n2366_o[18]\ _04549_ VPWR VGND _05776_ sg13g2_nor2_1
X_25506_ _04553_ _02045_ VPWR VGND _05777_ sg13g2_nor2_1
X_25507_ _02067_ _04533_ VPWR VGND _05778_ sg13g2_nor2_1
X_25508_ _04531_ _05777_ _05778_ _04536_ VPWR VGND 
+ _05779_
+ sg13g2_a22oi_1
X_25509_ _02045_ _04559_ VPWR VGND _05780_ sg13g2_nand2b_1
X_25510_ _04539_ _02067_ _05780_ VPWR VGND _05781_ sg13g2_o21ai_1
X_25511_ _04538_ _05781_ _04562_ VPWR VGND _05782_ sg13g2_a21oi_1
X_25512_ _04530_ _05779_ _05782_ VPWR VGND _05783_ sg13g2_a21oi_1
X_25513_ _04604_ _05775_ _05776_ _05783_ VPWR VGND 
+ _05784_
+ sg13g2_nor4_1
X_25514_ _04504_ _05774_ _05784_ VPWR VGND _05785_ sg13g2_nor3_1
X_25515_ \atbs_core_0.spike_memory_0.n2365_o[18]\ _04506_ VPWR VGND _05786_ sg13g2_nor2_1
X_25516_ \atbs_core_0.spike_memory_0.n2362_o[18]\ _04549_ VPWR VGND _05787_ sg13g2_nor2_1
X_25517_ _04553_ _12621_ VPWR VGND _05788_ sg13g2_nor2_1
X_25518_ _02019_ _04555_ VPWR VGND _05789_ sg13g2_nor2_1
X_25519_ _04378_ _05788_ _05789_ _04557_ VPWR VGND 
+ _05790_
+ sg13g2_a22oi_1
X_25520_ _12621_ _05544_ VPWR VGND _05791_ sg13g2_nand2b_1
X_25521_ _03755_ _02019_ _05791_ VPWR VGND _05792_ sg13g2_o21ai_1
X_25522_ _04388_ _05792_ _04562_ VPWR VGND _05793_ sg13g2_a21oi_1
X_25523_ _04551_ _05790_ _05793_ VPWR VGND _05794_ sg13g2_a21oi_1
X_25524_ _03729_ _05786_ _05787_ _05794_ VPWR VGND 
+ _05795_
+ sg13g2_nor4_1
X_25525_ \atbs_core_0.spike_memory_0.n2373_o[18]\ _12088_ VPWR VGND _05796_ sg13g2_nor2_1
X_25526_ \atbs_core_0.spike_memory_0.n2370_o[18]\ _04528_ VPWR VGND _05797_ sg13g2_nor2_1
X_25527_ _03934_ _02101_ VPWR VGND _05798_ sg13g2_nor2_1
X_25528_ _02124_ _04570_ VPWR VGND _05799_ sg13g2_nor2_1
X_25529_ _04568_ _05798_ _05799_ _02714_ VPWR VGND 
+ _05800_
+ sg13g2_a22oi_1
X_25530_ _02101_ _04361_ VPWR VGND _05801_ sg13g2_nand2b_1
X_25531_ _04574_ _02124_ _05801_ VPWR VGND _05802_ sg13g2_o21ai_1
X_25532_ _04573_ _05802_ _04338_ VPWR VGND _05803_ sg13g2_a21oi_1
X_25533_ _02702_ _05800_ _05803_ VPWR VGND _05804_ sg13g2_a21oi_1
X_25534_ _04126_ _05796_ _05797_ _05804_ VPWR VGND 
+ _05805_
+ sg13g2_nor4_1
X_25535_ _04547_ _05795_ _05805_ VPWR VGND _05806_ sg13g2_nor3_1
X_25536_ _07549_ _05785_ _05806_ VPWR VGND _05807_ sg13g2_nor3_1
X_25537_ _04333_ _05764_ _05807_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[18]\ sg13g2_a21o_1
X_25538_ _03754_ _02135_ VPWR VGND _05808_ sg13g2_nor2_1
X_25539_ _02158_ _03751_ VPWR VGND _05809_ sg13g2_nor2_1
X_25540_ _03744_ _05808_ _05809_ _04379_ VPWR VGND 
+ _05810_
+ sg13g2_a22oi_1
X_25541_ _02135_ _04111_ VPWR VGND _05811_ sg13g2_nand2b_1
X_25542_ _04512_ _02158_ _05811_ VPWR VGND _05812_ sg13g2_o21ai_1
X_25543_ _04387_ _05812_ _04392_ VPWR VGND _05813_ sg13g2_a21oi_1
X_25544_ _04376_ _05810_ _05813_ VPWR VGND _05814_ sg13g2_a21oi_1
X_25545_ _00115_ _03733_ _03737_ _02184_ _05814_ VPWR 
+ VGND
+ _05815_ sg13g2_a221oi_1
X_25546_ \atbs_core_0.spike_memory_0.n2385_o[1]\ _12086_ VPWR VGND _05816_ sg13g2_nor2_1
X_25547_ \atbs_core_0.spike_memory_0.n2382_o[1]\ _04771_ _03780_ VPWR VGND _05817_ sg13g2_o21ai_1
X_25548_ _03787_ _02287_ VPWR VGND _05818_ sg13g2_nor2_1
X_25549_ _02310_ _03785_ VPWR VGND _05819_ sg13g2_nor2_1
X_25550_ _03743_ _05818_ _05819_ _03754_ VPWR VGND 
+ _05820_
+ sg13g2_a22oi_1
X_25551_ _02287_ _03891_ VPWR VGND _05821_ sg13g2_nand2b_1
X_25552_ _03753_ _02310_ _05821_ VPWR VGND _05822_ sg13g2_o21ai_1
X_25553_ _03758_ _05822_ _04294_ VPWR VGND _05823_ sg13g2_a21oi_1
X_25554_ _03739_ _05820_ _05823_ VPWR VGND _05824_ sg13g2_a21oi_1
X_25555_ _05816_ _05817_ _05824_ VPWR VGND _05825_ sg13g2_or3_1
X_25556_ _03775_ _05825_ VPWR VGND _05826_ sg13g2_nand2_1
X_25557_ _03729_ _05815_ _05826_ VPWR VGND _05827_ sg13g2_o21ai_1
X_25558_ \atbs_core_0.spike_memory_0.n2381_o[1]\ _03944_ VPWR VGND _05828_ sg13g2_nor2_1
X_25559_ \atbs_core_0.spike_memory_0.n2378_o[1]\ _03807_ VPWR VGND _05829_ sg13g2_nor2_1
X_25560_ _03822_ _02233_ VPWR VGND _05830_ sg13g2_nor2_1
X_25561_ _02255_ _03909_ VPWR VGND _05831_ sg13g2_nor2_1
X_25562_ _04150_ _05830_ _05831_ _04154_ VPWR VGND 
+ _05832_
+ sg13g2_a22oi_1
X_25563_ _02233_ _05745_ VPWR VGND _05833_ sg13g2_nand2b_1
X_25564_ _05753_ _02255_ _05833_ VPWR VGND _05834_ sg13g2_o21ai_1
X_25565_ _03913_ _05834_ _03919_ VPWR VGND _05835_ sg13g2_a21oi_1
X_25566_ _04149_ _05832_ _05835_ VPWR VGND _05836_ sg13g2_a21oi_1
X_25567_ _05828_ _05829_ _05836_ VPWR VGND _05837_ sg13g2_nor3_1
X_25568_ \atbs_core_0.spike_memory_0.n2389_o[1]\ _03736_ VPWR VGND _05838_ sg13g2_nand2b_1
X_25569_ \atbs_core_0.spike_memory_0.n2386_o[1]\ _03836_ _05838_ VPWR VGND _05839_ sg13g2_o21ai_1
X_25570_ _03856_ _02343_ VPWR VGND _05840_ sg13g2_nor2_1
X_25571_ _02367_ _03952_ VPWR VGND _05841_ sg13g2_nor2_1
X_25572_ _03844_ _05840_ _05841_ _03857_ VPWR VGND 
+ _05842_
+ sg13g2_a22oi_1
X_25573_ _02343_ _04167_ VPWR VGND _05843_ sg13g2_nand2b_1
X_25574_ _03949_ _02367_ _05843_ VPWR VGND _05844_ sg13g2_o21ai_1
X_25575_ _03956_ _05844_ _04317_ VPWR VGND _05845_ sg13g2_a21oi_1
X_25576_ _03841_ _05842_ _05845_ VPWR VGND _05846_ sg13g2_a21oi_1
X_25577_ _05839_ _05846_ _03775_ VPWR VGND _05847_ sg13g2_o21ai_1
X_25578_ _03801_ _05837_ _05847_ VPWR VGND _05848_ sg13g2_o21ai_1
X_25579_ _03725_ _05827_ _05848_ _05825_ VPWR VGND 
+ _05849_
+ sg13g2_a22oi_1
X_25580_ _04254_ VPWR VGND _05850_ sg13g2_buf_1
X_25581_ _05850_ _02619_ VPWR VGND _05851_ sg13g2_nor2_1
X_25582_ _02640_ _04047_ VPWR VGND _05852_ sg13g2_nor2_1
X_25583_ _04587_ _05851_ _05852_ _04610_ VPWR VGND 
+ _05853_
+ sg13g2_a22oi_1
X_25584_ _02619_ _05533_ VPWR VGND _05854_ sg13g2_nand2b_1
X_25585_ _03983_ _02640_ _05854_ VPWR VGND _05855_ sg13g2_o21ai_1
X_25586_ _03987_ _05855_ _03811_ VPWR VGND _05856_ sg13g2_a21oi_1
X_25587_ _03974_ _05853_ _05856_ VPWR VGND _05857_ sg13g2_a21oi_1
X_25588_ _00113_ _03969_ _03972_ _02662_ _05857_ VPWR 
+ VGND
+ _05858_ sg13g2_a221oi_1
X_25589_ \atbs_core_0.spike_memory_0.n2417_o[1]\ _03876_ VPWR VGND _05859_ sg13g2_nor2_1
X_25590_ \atbs_core_0.spike_memory_0.n2414_o[1]\ _04229_ _03722_ VPWR VGND _05860_ sg13g2_o21ai_1
X_25591_ _03977_ _12573_ VPWR VGND _05861_ sg13g2_nor2_1
X_25592_ _12596_ _04062_ VPWR VGND _05862_ sg13g2_nor2_1
X_25593_ _03975_ _05861_ _05862_ _05850_ VPWR VGND 
+ _05863_
+ sg13g2_a22oi_1
X_25594_ _12573_ _04088_ VPWR VGND _05864_ sg13g2_nand2b_1
X_25595_ _04094_ _12596_ _05864_ VPWR VGND _05865_ sg13g2_o21ai_1
X_25596_ _04010_ _05865_ _03992_ VPWR VGND _05866_ sg13g2_a21oi_1
X_25597_ _04002_ _05863_ _05866_ VPWR VGND _05867_ sg13g2_a21oi_1
X_25598_ _05859_ _05860_ _05867_ VPWR VGND _05868_ sg13g2_or3_1
X_25599_ _03926_ _05868_ VPWR VGND _05869_ sg13g2_nand2_1
X_25600_ _03968_ _05858_ _05869_ VPWR VGND _05870_ sg13g2_o21ai_1
X_25601_ \atbs_core_0.spike_memory_0.n2413_o[1]\ _12087_ VPWR VGND _05871_ sg13g2_nor2_1
X_25602_ \atbs_core_0.spike_memory_0.n2410_o[1]\ _04527_ VPWR VGND _05872_ sg13g2_nor2_1
X_25603_ _03886_ _12517_ VPWR VGND _05873_ sg13g2_nor2_1
X_25604_ _12541_ _04082_ VPWR VGND _05874_ sg13g2_nor2_1
X_25605_ _04359_ _05873_ _05874_ _04535_ VPWR VGND 
+ _05875_
+ sg13g2_a22oi_1
X_25606_ _12517_ _04105_ VPWR VGND _05876_ sg13g2_nand2b_1
X_25607_ _03747_ _12541_ _05876_ VPWR VGND _05877_ sg13g2_o21ai_1
X_25608_ _03759_ _05877_ _03769_ VPWR VGND _05878_ sg13g2_a21oi_1
X_25609_ _03740_ _05875_ _05878_ VPWR VGND _05879_ sg13g2_a21oi_1
X_25610_ _05871_ _05872_ _05879_ VPWR VGND _05880_ sg13g2_nor3_1
X_25611_ \atbs_core_0.spike_memory_0.n2436_q[1198]\ _03971_ VPWR VGND _05881_ sg13g2_nand2b_1
X_25612_ \atbs_core_0.spike_memory_0.n2418_o[1]\ _04032_ _05881_ VPWR VGND _05882_ sg13g2_o21ai_1
X_25613_ _03826_ _12631_ VPWR VGND _05883_ sg13g2_nor2_1
X_25614_ _12654_ _03932_ VPWR VGND _05884_ sg13g2_nor2_1
X_25615_ _03929_ _05883_ _05884_ _04154_ VPWR VGND 
+ _05885_
+ sg13g2_a22oi_1
X_25616_ _12631_ _03937_ VPWR VGND _05886_ sg13g2_nand2b_1
X_25617_ _02712_ _12654_ _05886_ VPWR VGND _05887_ sg13g2_o21ai_1
X_25618_ _03936_ _05887_ _04158_ VPWR VGND _05888_ sg13g2_a21oi_1
X_25619_ _02701_ _05885_ _05888_ VPWR VGND _05889_ sg13g2_a21oi_1
X_25620_ _05882_ _05889_ _03997_ VPWR VGND _05890_ sg13g2_o21ai_1
X_25621_ _03801_ _05880_ _05890_ VPWR VGND _05891_ sg13g2_o21ai_1
X_25622_ _03967_ _05870_ _05891_ _05868_ _04045_ VPWR 
+ VGND
+ _05892_ sg13g2_a221oi_1
X_25623_ _03721_ _05849_ _05892_ VPWR VGND _05893_ sg13g2_a21oi_1
X_25624_ \atbs_core_0.spike_memory_0.n2369_o[1]\ _03803_ VPWR VGND _05894_ sg13g2_nor2_1
X_25625_ \atbs_core_0.spike_memory_0.n2366_o[1]\ _03806_ VPWR VGND _05895_ sg13g2_nor2_1
X_25626_ _03815_ _02025_ VPWR VGND _05896_ sg13g2_nor2_1
X_25627_ _02048_ _03951_ VPWR VGND _05897_ sg13g2_nor2_1
X_25628_ _03813_ _05896_ _05897_ _03907_ VPWR VGND 
+ _05898_
+ sg13g2_a22oi_1
X_25629_ _02025_ _03915_ VPWR VGND _05899_ sg13g2_nand2b_1
X_25630_ _03821_ _02048_ _05899_ VPWR VGND _05900_ sg13g2_o21ai_1
X_25631_ _03790_ _05900_ _03830_ VPWR VGND _05901_ sg13g2_a21oi_1
X_25632_ _03811_ _05898_ _05901_ VPWR VGND _05902_ sg13g2_a21oi_1
X_25633_ _05894_ _05895_ _05902_ VPWR VGND _05903_ sg13g2_nor3_1
X_25634_ \atbs_core_0.spike_memory_0.n2361_o[1]\ _03803_ VPWR VGND _05904_ sg13g2_nor2_1
X_25635_ \atbs_core_0.spike_memory_0.n2358_o[1]\ _05540_ VPWR VGND _05905_ sg13g2_nor2_1
X_25636_ _03855_ _02069_ VPWR VGND _05906_ sg13g2_nor2_1
X_25637_ _02232_ _03851_ VPWR VGND _05907_ sg13g2_nor2_1
X_25638_ _03843_ _05906_ _05907_ _03949_ VPWR VGND 
+ _05908_
+ sg13g2_a22oi_1
X_25639_ _02069_ _04054_ VPWR VGND _05909_ sg13g2_nand2b_1
X_25640_ _04051_ _02232_ _05909_ VPWR VGND _05910_ sg13g2_o21ai_1
X_25641_ _03955_ _05910_ _03868_ VPWR VGND _05911_ sg13g2_a21oi_1
X_25642_ _03993_ _05908_ _05911_ VPWR VGND _05912_ sg13g2_a21oi_1
X_25643_ _04244_ _05904_ _05905_ _05912_ VPWR VGND 
+ _05913_
+ sg13g2_nor4_1
X_25644_ _03926_ _05903_ _05913_ VPWR VGND _05914_ sg13g2_a21oi_1
X_25645_ \atbs_core_0.spike_memory_0.n2365_o[1]\ _03776_ VPWR VGND _05915_ sg13g2_nor2_1
X_25646_ \atbs_core_0.spike_memory_0.n2362_o[1]\ _03806_ VPWR VGND _05916_ sg13g2_nor2_1
X_25647_ _03855_ _12630_ VPWR VGND _05917_ sg13g2_nor2_1
X_25648_ _12629_ _03951_ VPWR VGND _05918_ sg13g2_nor2_1
X_25649_ _04047_ _05917_ _05918_ _03957_ VPWR VGND 
+ _05919_
+ sg13g2_a22oi_1
X_25650_ _12630_ _04054_ VPWR VGND _05920_ sg13g2_nand2b_1
X_25651_ _03815_ _12629_ _05920_ VPWR VGND _05921_ sg13g2_o21ai_1
X_25652_ _03955_ _05921_ _03868_ VPWR VGND _05922_ sg13g2_a21oi_1
X_25653_ _03993_ _05919_ _05922_ VPWR VGND _05923_ sg13g2_a21oi_1
X_25654_ _04244_ _05915_ _05916_ _05923_ VPWR VGND 
+ _05924_
+ sg13g2_nor4_1
X_25655_ \atbs_core_0.spike_memory_0.n2373_o[1]\ _03803_ VPWR VGND _05925_ sg13g2_nor2_1
X_25656_ \atbs_core_0.spike_memory_0.n2370_o[1]\ _04102_ VPWR VGND _05926_ sg13g2_nor2_1
X_25657_ _05533_ _02080_ VPWR VGND _05927_ sg13g2_nor2_1
X_25658_ _02103_ _03851_ VPWR VGND _05928_ sg13g2_nor2_1
X_25659_ _03843_ _05927_ _05928_ _04708_ VPWR VGND 
+ _05929_
+ sg13g2_a22oi_1
X_25660_ _02080_ _03982_ VPWR VGND _05930_ sg13g2_nand2b_1
X_25661_ _04597_ _02103_ _05930_ VPWR VGND _05931_ sg13g2_o21ai_1
X_25662_ _03860_ _05931_ _04287_ VPWR VGND _05932_ sg13g2_a21oi_1
X_25663_ _03840_ _05929_ _05932_ VPWR VGND _05933_ sg13g2_a21oi_1
X_25664_ _03899_ _05925_ _05926_ _05933_ VPWR VGND 
+ _05934_
+ sg13g2_nor4_1
X_25665_ _03724_ _05924_ _05934_ VPWR VGND _05935_ sg13g2_nor3_1
X_25666_ _03724_ _05914_ _05935_ VPWR VGND _05936_ sg13g2_a21oi_1
X_25667_ _04045_ _05936_ VPWR VGND _05937_ sg13g2_and2_1
X_25668_ _05850_ _02392_ VPWR VGND _05938_ sg13g2_nor2_1
X_25669_ _02412_ _04047_ VPWR VGND _05939_ sg13g2_nor2_1
X_25670_ _04587_ _05938_ _05939_ _03984_ VPWR VGND 
+ _05940_
+ sg13g2_a22oi_1
X_25671_ _02392_ _03989_ VPWR VGND _05941_ sg13g2_nand2b_1
X_25672_ _03983_ _02412_ _05941_ VPWR VGND _05942_ sg13g2_o21ai_1
X_25673_ _03987_ _05942_ _03811_ VPWR VGND _05943_ sg13g2_a21oi_1
X_25674_ _03974_ _05940_ _05943_ VPWR VGND _05944_ sg13g2_a21oi_1
X_25675_ _00114_ _03969_ _03972_ _02432_ _05944_ VPWR 
+ VGND
+ _05945_ sg13g2_a221oi_1
X_25676_ \atbs_core_0.spike_memory_0.n2401_o[1]\ _03876_ VPWR VGND _05946_ sg13g2_nor2_1
X_25677_ \atbs_core_0.spike_memory_0.n2398_o[1]\ _04229_ _03722_ VPWR VGND _05947_ sg13g2_o21ai_1
X_25678_ _03977_ _02524_ VPWR VGND _05948_ sg13g2_nor2_1
X_25679_ _02545_ _04062_ VPWR VGND _05949_ sg13g2_nor2_1
X_25680_ _03975_ _05948_ _05949_ _05850_ VPWR VGND 
+ _05950_
+ sg13g2_a22oi_1
X_25681_ _02524_ _04011_ VPWR VGND _05951_ sg13g2_nand2b_1
X_25682_ _04254_ _02545_ _05951_ VPWR VGND _05952_ sg13g2_o21ai_1
X_25683_ _04010_ _05952_ _03839_ VPWR VGND _05953_ sg13g2_a21oi_1
X_25684_ _04002_ _05950_ _05953_ VPWR VGND _05954_ sg13g2_a21oi_1
X_25685_ _05946_ _05947_ _05954_ VPWR VGND _05955_ sg13g2_or3_1
X_25686_ _03997_ _05955_ VPWR VGND _05956_ sg13g2_nand2_1
X_25687_ _03968_ _05945_ _05956_ VPWR VGND _05957_ sg13g2_o21ai_1
X_25688_ \atbs_core_0.spike_memory_0.n2397_o[1]\ _12087_ VPWR VGND _05958_ sg13g2_nor2_1
X_25689_ \atbs_core_0.spike_memory_0.n2394_o[1]\ _03836_ VPWR VGND _05959_ sg13g2_nor2_1
X_25690_ _04552_ _02476_ VPWR VGND _05960_ sg13g2_nor2_1
X_25691_ _02498_ _04023_ VPWR VGND _05961_ sg13g2_nor2_1
X_25692_ _04359_ _05960_ _05961_ _04535_ VPWR VGND 
+ _05962_
+ sg13g2_a22oi_1
X_25693_ _02476_ _04105_ VPWR VGND _05963_ sg13g2_nand2b_1
X_25694_ _03788_ _02498_ _05963_ VPWR VGND _05964_ sg13g2_o21ai_1
X_25695_ _03759_ _05964_ _04081_ VPWR VGND _05965_ sg13g2_a21oi_1
X_25696_ _04021_ _05962_ _05965_ VPWR VGND _05966_ sg13g2_a21oi_1
X_25697_ _05958_ _05959_ _05966_ VPWR VGND _05967_ sg13g2_nor3_1
X_25698_ \atbs_core_0.spike_memory_0.n2405_o[1]\ _03971_ VPWR VGND _05968_ sg13g2_nand2b_1
X_25699_ \atbs_core_0.spike_memory_0.n2402_o[1]\ _04032_ _05968_ VPWR VGND _05969_ sg13g2_o21ai_1
X_25700_ _03826_ _02572_ VPWR VGND _05970_ sg13g2_nor2_1
X_25701_ _02593_ _04152_ VPWR VGND _05971_ sg13g2_nor2_1
X_25702_ _04150_ _05970_ _05971_ _04154_ VPWR VGND 
+ _05972_
+ sg13g2_a22oi_1
X_25703_ _02572_ _05745_ VPWR VGND _05973_ sg13g2_nand2b_1
X_25704_ _05753_ _02593_ _05973_ VPWR VGND _05974_ sg13g2_o21ai_1
X_25705_ _03936_ _05974_ _04158_ VPWR VGND _05975_ sg13g2_a21oi_1
X_25706_ _04149_ _05972_ _05975_ VPWR VGND _05976_ sg13g2_a21oi_1
X_25707_ _05969_ _05976_ _03997_ VPWR VGND _05977_ sg13g2_o21ai_1
X_25708_ _03801_ _05967_ _05977_ VPWR VGND _05978_ sg13g2_o21ai_1
X_25709_ _03967_ _05957_ _05978_ _05955_ _04045_ VPWR 
+ VGND
+ _05979_ sg13g2_a221oi_1
X_25710_ _05937_ _05979_ _03719_ VPWR VGND _05980_ sg13g2_o21ai_1
X_25711_ _03719_ _05893_ _05980_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[1]\ sg13g2_o21ai_1
X_25712_ _03761_ _02136_ VPWR VGND _05981_ sg13g2_nor2_1
X_25713_ _02160_ _03751_ VPWR VGND _05982_ sg13g2_nor2_1
X_25714_ _03744_ _05981_ _05982_ _04379_ VPWR VGND 
+ _05983_
+ sg13g2_a22oi_1
X_25715_ _02136_ _04111_ VPWR VGND _05984_ sg13g2_nand2b_1
X_25716_ _04512_ _02160_ _05984_ VPWR VGND _05985_ sg13g2_o21ai_1
X_25717_ _04387_ _05985_ _03840_ VPWR VGND _05986_ sg13g2_a21oi_1
X_25718_ _04376_ _05983_ _05986_ VPWR VGND _05987_ sg13g2_a21oi_1
X_25719_ _00118_ _03733_ _03737_ _02186_ _05987_ VPWR 
+ VGND
+ _05988_ sg13g2_a221oi_1
X_25720_ \atbs_core_0.spike_memory_0.n2385_o[2]\ _12086_ VPWR VGND _05989_ sg13g2_nor2_1
X_25721_ \atbs_core_0.spike_memory_0.n2382_o[2]\ _04771_ _03780_ VPWR VGND _05990_ sg13g2_o21ai_1
X_25722_ _03787_ _02288_ VPWR VGND _05991_ sg13g2_nor2_1
X_25723_ _02311_ _03750_ VPWR VGND _05992_ sg13g2_nor2_1
X_25724_ _03743_ _05991_ _05992_ _03754_ VPWR VGND 
+ _05993_
+ sg13g2_a22oi_1
X_25725_ _02288_ _03763_ VPWR VGND _05994_ sg13g2_nand2b_1
X_25726_ _03753_ _02311_ _05994_ VPWR VGND _05995_ sg13g2_o21ai_1
X_25727_ _03758_ _05995_ _04294_ VPWR VGND _05996_ sg13g2_a21oi_1
X_25728_ _03739_ _05993_ _05996_ VPWR VGND _05997_ sg13g2_a21oi_1
X_25729_ _05989_ _05990_ _05997_ VPWR VGND _05998_ sg13g2_or3_1
X_25730_ _03775_ _05998_ VPWR VGND _05999_ sg13g2_nand2_1
X_25731_ _03729_ _05988_ _05999_ VPWR VGND _06000_ sg13g2_o21ai_1
X_25732_ \atbs_core_0.spike_memory_0.n2381_o[2]\ _03944_ VPWR VGND _06001_ sg13g2_nor2_1
X_25733_ \atbs_core_0.spike_memory_0.n2378_o[2]\ _03807_ VPWR VGND _06002_ sg13g2_nor2_1
X_25734_ _03822_ _02234_ VPWR VGND _06003_ sg13g2_nor2_1
X_25735_ _02257_ _04152_ VPWR VGND _06004_ sg13g2_nor2_1
X_25736_ _04150_ _06003_ _06004_ _04154_ VPWR VGND 
+ _06005_
+ sg13g2_a22oi_1
X_25737_ _02234_ _05745_ VPWR VGND _06006_ sg13g2_nand2b_1
X_25738_ _05753_ _02257_ _06006_ VPWR VGND _06007_ sg13g2_o21ai_1
X_25739_ _03936_ _06007_ _04158_ VPWR VGND _06008_ sg13g2_a21oi_1
X_25740_ _04149_ _06005_ _06008_ VPWR VGND _06009_ sg13g2_a21oi_1
X_25741_ _06001_ _06002_ _06009_ VPWR VGND _06010_ sg13g2_nor3_1
X_25742_ \atbs_core_0.spike_memory_0.n2389_o[2]\ _03971_ VPWR VGND _06011_ sg13g2_nand2b_1
X_25743_ \atbs_core_0.spike_memory_0.n2386_o[2]\ _03836_ _06011_ VPWR VGND _06012_ sg13g2_o21ai_1
X_25744_ _03856_ _02344_ VPWR VGND _06013_ sg13g2_nor2_1
X_25745_ _02368_ _03952_ VPWR VGND _06014_ sg13g2_nor2_1
X_25746_ _03844_ _06013_ _06014_ _03857_ VPWR VGND 
+ _06015_
+ sg13g2_a22oi_1
X_25747_ _02344_ _04167_ VPWR VGND _06016_ sg13g2_nand2b_1
X_25748_ _03949_ _02368_ _06016_ VPWR VGND _06017_ sg13g2_o21ai_1
X_25749_ _03956_ _06017_ _04317_ VPWR VGND _06018_ sg13g2_a21oi_1
X_25750_ _03841_ _06015_ _06018_ VPWR VGND _06019_ sg13g2_a21oi_1
X_25751_ _06012_ _06019_ _03775_ VPWR VGND _06020_ sg13g2_o21ai_1
X_25752_ _03801_ _06010_ _06020_ VPWR VGND _06021_ sg13g2_o21ai_1
X_25753_ _03725_ _06000_ _06021_ _05998_ VPWR VGND 
+ _06022_
+ sg13g2_a22oi_1
X_25754_ _05850_ _02620_ VPWR VGND _06023_ sg13g2_nor2_1
X_25755_ _02641_ _04047_ VPWR VGND _06024_ sg13g2_nor2_1
X_25756_ _04587_ _06023_ _06024_ _04610_ VPWR VGND 
+ _06025_
+ sg13g2_a22oi_1
X_25757_ _02620_ _05533_ VPWR VGND _06026_ sg13g2_nand2b_1
X_25758_ _04589_ _02641_ _06026_ VPWR VGND _06027_ sg13g2_o21ai_1
X_25759_ _03987_ _06027_ _03811_ VPWR VGND _06028_ sg13g2_a21oi_1
X_25760_ _03974_ _06025_ _06028_ VPWR VGND _06029_ sg13g2_a21oi_1
X_25761_ _00116_ _03969_ _03972_ _02664_ _06029_ VPWR 
+ VGND
+ _06030_ sg13g2_a221oi_1
X_25762_ \atbs_core_0.spike_memory_0.n2417_o[2]\ _03876_ VPWR VGND _06031_ sg13g2_nor2_1
X_25763_ \atbs_core_0.spike_memory_0.n2414_o[2]\ _04229_ _03722_ VPWR VGND _06032_ sg13g2_o21ai_1
X_25764_ _03977_ _12574_ VPWR VGND _06033_ sg13g2_nor2_1
X_25765_ _12597_ _04062_ VPWR VGND _06034_ sg13g2_nor2_1
X_25766_ _03975_ _06033_ _06034_ _05850_ VPWR VGND 
+ _06035_
+ sg13g2_a22oi_1
X_25767_ _12574_ _04088_ VPWR VGND _06036_ sg13g2_nand2b_1
X_25768_ _04094_ _12597_ _06036_ VPWR VGND _06037_ sg13g2_o21ai_1
X_25769_ _04010_ _06037_ _03992_ VPWR VGND _06038_ sg13g2_a21oi_1
X_25770_ _04002_ _06035_ _06038_ VPWR VGND _06039_ sg13g2_a21oi_1
X_25771_ _06031_ _06032_ _06039_ VPWR VGND _06040_ sg13g2_or3_1
X_25772_ _03926_ _06040_ VPWR VGND _06041_ sg13g2_nand2_1
X_25773_ _03968_ _06030_ _06041_ VPWR VGND _06042_ sg13g2_o21ai_1
X_25774_ \atbs_core_0.spike_memory_0.n2413_o[2]\ _03877_ VPWR VGND _06043_ sg13g2_nor2_1
X_25775_ \atbs_core_0.spike_memory_0.n2410_o[2]\ _04527_ VPWR VGND _06044_ sg13g2_nor2_1
X_25776_ _03886_ _12518_ VPWR VGND _06045_ sg13g2_nor2_1
X_25777_ _12542_ _04082_ VPWR VGND _06046_ sg13g2_nor2_1
X_25778_ _04359_ _06045_ _06046_ _04535_ VPWR VGND 
+ _06047_
+ sg13g2_a22oi_1
X_25779_ _12518_ _04105_ VPWR VGND _06048_ sg13g2_nand2b_1
X_25780_ _03747_ _12542_ _06048_ VPWR VGND _06049_ sg13g2_o21ai_1
X_25781_ _03759_ _06049_ _03769_ VPWR VGND _06050_ sg13g2_a21oi_1
X_25782_ _03740_ _06047_ _06050_ VPWR VGND _06051_ sg13g2_a21oi_1
X_25783_ _06043_ _06044_ _06051_ VPWR VGND _06052_ sg13g2_nor3_1
X_25784_ \atbs_core_0.spike_memory_0.n2436_q[1199]\ _03971_ VPWR VGND _06053_ sg13g2_nand2b_1
X_25785_ \atbs_core_0.spike_memory_0.n2418_o[2]\ _04032_ _06053_ VPWR VGND _06054_ sg13g2_o21ai_1
X_25786_ _03826_ _12632_ VPWR VGND _06055_ sg13g2_nor2_1
X_25787_ _12657_ _03932_ VPWR VGND _06056_ sg13g2_nor2_1
X_25788_ _03929_ _06055_ _06056_ _04154_ VPWR VGND 
+ _06057_
+ sg13g2_a22oi_1
X_25789_ _12632_ _03937_ VPWR VGND _06058_ sg13g2_nand2b_1
X_25790_ _02712_ _12657_ _06058_ VPWR VGND _06059_ sg13g2_o21ai_1
X_25791_ _03936_ _06059_ _04158_ VPWR VGND _06060_ sg13g2_a21oi_1
X_25792_ _02701_ _06057_ _06060_ VPWR VGND _06061_ sg13g2_a21oi_1
X_25793_ _06054_ _06061_ _03997_ VPWR VGND _06062_ sg13g2_o21ai_1
X_25794_ _04074_ _06052_ _06062_ VPWR VGND _06063_ sg13g2_o21ai_1
X_25795_ _03967_ _06042_ _06063_ _06040_ _04045_ VPWR 
+ VGND
+ _06064_ sg13g2_a221oi_1
X_25796_ _03721_ _06022_ _06064_ VPWR VGND _06065_ sg13g2_a21oi_1
X_25797_ \atbs_core_0.spike_memory_0.n2392_o[2]\ _03986_ VPWR VGND _06066_ sg13g2_nand2_1
X_25798_ _00117_ _03860_ _06066_ VPWR VGND _06067_ sg13g2_o21ai_1
X_25799_ _07528_ _07560_ _04003_ VPWR VGND _06068_ sg13g2_mux2_1
X_25800_ _07561_ _06067_ _06068_ \atbs_core_0.spike_memory_0.n2391_o[2]\ VPWR VGND 
+ _06069_
+ sg13g2_a22oi_1
X_25801_ _02435_ _03804_ _06069_ VPWR VGND _06070_ sg13g2_o21ai_1
X_25802_ \atbs_core_0.spike_memory_0.n2401_o[2]\ _04260_ VPWR VGND _06071_ sg13g2_nor2_1
X_25803_ \atbs_core_0.spike_memory_0.n2398_o[2]\ _04230_ VPWR VGND _06072_ sg13g2_nor2_1
X_25804_ _04346_ _02525_ VPWR VGND _06073_ sg13g2_nor2_1
X_25805_ _02546_ _04265_ VPWR VGND _06074_ sg13g2_nor2_1
X_25806_ _05496_ _06073_ _06074_ _04112_ VPWR VGND 
+ _06075_
+ sg13g2_a22oi_1
X_25807_ _02525_ _03760_ VPWR VGND _06076_ sg13g2_nand2b_1
X_25808_ _04236_ _02546_ _06076_ VPWR VGND _06077_ sg13g2_o21ai_1
X_25809_ _04235_ _06077_ _03973_ VPWR VGND _06078_ sg13g2_a21oi_1
X_25810_ _03940_ _06075_ _06078_ VPWR VGND _06079_ sg13g2_a21oi_1
X_25811_ _03899_ _06071_ _06072_ _06079_ VPWR VGND 
+ _06080_
+ sg13g2_nor4_1
X_25812_ _04219_ _06070_ _06080_ VPWR VGND _06081_ sg13g2_a21oi_1
X_25813_ \atbs_core_0.spike_memory_0.n2397_o[2]\ _04245_ VPWR VGND _06082_ sg13g2_nor2_1
X_25814_ \atbs_core_0.spike_memory_0.n2394_o[2]\ _04247_ VPWR VGND _06083_ sg13g2_nor2_1
X_25815_ _04083_ _02477_ VPWR VGND _06084_ sg13g2_nor2_1
X_25816_ _02499_ _04250_ VPWR VGND _06085_ sg13g2_nor2_1
X_25817_ _04082_ _06084_ _06085_ _04090_ VPWR VGND 
+ _06086_
+ sg13g2_a22oi_1
X_25818_ _02477_ _04254_ VPWR VGND _06087_ sg13g2_nand2b_1
X_25819_ _04089_ _02499_ _06087_ VPWR VGND _06088_ sg13g2_o21ai_1
X_25820_ _04253_ _06088_ _04098_ VPWR VGND _06089_ sg13g2_a21oi_1
X_25821_ _04081_ _06086_ _06089_ VPWR VGND _06090_ sg13g2_a21oi_1
X_25822_ _04244_ _06082_ _06083_ _06090_ VPWR VGND 
+ _06091_
+ sg13g2_nor4_1
X_25823_ \atbs_core_0.spike_memory_0.n2405_o[2]\ _04260_ VPWR VGND _06092_ sg13g2_nor2_1
X_25824_ \atbs_core_0.spike_memory_0.n2402_o[2]\ _04079_ VPWR VGND _06093_ sg13g2_nor2_1
X_25825_ _04236_ _02573_ VPWR VGND _06094_ sg13g2_nor2_1
X_25826_ _02594_ _04250_ VPWR VGND _06095_ sg13g2_nor2_1
X_25827_ _03884_ _06094_ _06095_ _04518_ VPWR VGND 
+ _06096_
+ sg13g2_a22oi_1
X_25828_ _02573_ _03977_ VPWR VGND _06097_ sg13g2_nand2b_1
X_25829_ _04083_ _02594_ _06097_ VPWR VGND _06098_ sg13g2_o21ai_1
X_25830_ _04253_ _06098_ _04272_ VPWR VGND _06099_ sg13g2_a21oi_1
X_25831_ _03895_ _06096_ _06099_ VPWR VGND _06100_ sg13g2_a21oi_1
X_25832_ _03899_ _06092_ _06093_ _06100_ VPWR VGND 
+ _06101_
+ sg13g2_nor4_1
X_25833_ _06091_ _06101_ _04277_ VPWR VGND _06102_ sg13g2_o21ai_1
X_25834_ _03925_ _06081_ _06102_ VPWR VGND _06103_ sg13g2_o21ai_1
X_25835_ \atbs_core_0.spike_memory_0.n2369_o[2]\ _04076_ VPWR VGND _06104_ sg13g2_nor2_1
X_25836_ \atbs_core_0.spike_memory_0.n2366_o[2]\ _04079_ VPWR VGND _06105_ sg13g2_nor2_1
X_25837_ _04267_ _02028_ VPWR VGND _06106_ sg13g2_nor2_1
X_25838_ _02049_ _04250_ VPWR VGND _06107_ sg13g2_nor2_1
X_25839_ _04023_ _06106_ _06107_ _04090_ VPWR VGND 
+ _06108_
+ sg13g2_a22oi_1
X_25840_ _02028_ _03977_ VPWR VGND _06109_ sg13g2_nand2b_1
X_25841_ _04089_ _02049_ _06109_ VPWR VGND _06110_ sg13g2_o21ai_1
X_25842_ _04253_ _06110_ _04272_ VPWR VGND _06111_ sg13g2_a21oi_1
X_25843_ _03895_ _06108_ _06111_ VPWR VGND _06112_ sg13g2_a21oi_1
X_25844_ _06104_ _06105_ _06112_ VPWR VGND _06113_ sg13g2_nor3_1
X_25845_ \atbs_core_0.spike_memory_0.n2361_o[2]\ _04076_ VPWR VGND _06114_ sg13g2_nor2_1
X_25846_ \atbs_core_0.spike_memory_0.n2358_o[2]\ _04230_ VPWR VGND _06115_ sg13g2_nor2_1
X_25847_ _04346_ _02071_ VPWR VGND _06116_ sg13g2_nor2_1
X_25848_ _02244_ _04108_ VPWR VGND _06117_ sg13g2_nor2_1
X_25849_ _03932_ _06116_ _06117_ _04112_ VPWR VGND 
+ _06118_
+ sg13g2_a22oi_1
X_25850_ _02071_ _04237_ VPWR VGND _06119_ sg13g2_nand2b_1
X_25851_ _04236_ _02244_ _06119_ VPWR VGND _06120_ sg13g2_o21ai_1
X_25852_ _04235_ _06120_ _03973_ VPWR VGND _06121_ sg13g2_a21oi_1
X_25853_ _03940_ _06118_ _06121_ VPWR VGND _06122_ sg13g2_a21oi_1
X_25854_ _03774_ _06114_ _06115_ _06122_ VPWR VGND 
+ _06123_
+ sg13g2_nor4_1
X_25855_ _03997_ _06113_ _06123_ VPWR VGND _06124_ sg13g2_a21oi_1
X_25856_ \atbs_core_0.spike_memory_0.n2365_o[2]\ _04260_ VPWR VGND _06125_ sg13g2_nor2_1
X_25857_ \atbs_core_0.spike_memory_0.n2362_o[2]\ _04079_ VPWR VGND _06126_ sg13g2_nor2_1
X_25858_ _04111_ _12643_ VPWR VGND _06127_ sg13g2_nor2_1
X_25859_ _12642_ _04265_ VPWR VGND _06128_ sg13g2_nor2_1
X_25860_ _03884_ _06127_ _06128_ _04268_ VPWR VGND 
+ _06129_
+ sg13g2_a22oi_1
X_25861_ _12643_ _04004_ VPWR VGND _06130_ sg13g2_nand2b_1
X_25862_ _04267_ _12642_ _06130_ VPWR VGND _06131_ sg13g2_o21ai_1
X_25863_ _04235_ _06131_ _04272_ VPWR VGND _06132_ sg13g2_a21oi_1
X_25864_ _04263_ _06129_ _06132_ VPWR VGND _06133_ sg13g2_a21oi_1
X_25865_ _03774_ _06125_ _06126_ _06133_ VPWR VGND 
+ _06134_
+ sg13g2_nor4_1
X_25866_ \atbs_core_0.spike_memory_0.n2373_o[2]\ _04076_ VPWR VGND _06135_ sg13g2_nor2_1
X_25867_ \atbs_core_0.spike_memory_0.n2370_o[2]\ _04230_ VPWR VGND _06136_ sg13g2_nor2_1
X_25868_ _03892_ _02081_ VPWR VGND _06137_ sg13g2_nor2_1
X_25869_ _02104_ _04003_ VPWR VGND _06138_ sg13g2_nor2_1
X_25870_ _03819_ _06137_ _06138_ _04347_ VPWR VGND 
+ _06139_
+ sg13g2_a22oi_1
X_25871_ _02081_ _03746_ VPWR VGND _06140_ sg13g2_nand2b_1
X_25872_ _04026_ _02104_ _06140_ VPWR VGND _06141_ sg13g2_o21ai_1
X_25873_ _04114_ _06141_ _04002_ VPWR VGND _06142_ sg13g2_a21oi_1
X_25874_ _03831_ _06139_ _06142_ VPWR VGND _06143_ sg13g2_a21oi_1
X_25875_ _03899_ _06135_ _06136_ _06143_ VPWR VGND 
+ _06144_
+ sg13g2_nor4_1
X_25876_ _03724_ _06134_ _06144_ VPWR VGND _06145_ sg13g2_nor3_1
X_25877_ _03967_ _06124_ _06145_ VPWR VGND _06146_ sg13g2_a21oi_1
X_25878_ _06103_ _06146_ _04330_ VPWR VGND _06147_ sg13g2_mux2_1
X_25879_ _03719_ _06147_ VPWR VGND _06148_ sg13g2_nand2_1
X_25880_ _03719_ _06065_ _06148_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[2]\ sg13g2_o21ai_1
X_25881_ _04340_ _02393_ VPWR VGND _06149_ sg13g2_nor2_1
X_25882_ _02413_ _03976_ VPWR VGND _06150_ sg13g2_nor2_1
X_25883_ _04339_ _06149_ _06150_ _04343_ VPWR VGND 
+ _06151_
+ sg13g2_a22oi_1
X_25884_ _02393_ _03788_ VPWR VGND _06152_ sg13g2_nand2b_1
X_25885_ _04347_ _02413_ _06152_ VPWR VGND _06153_ sg13g2_o21ai_1
X_25886_ _04345_ _06153_ _04684_ VPWR VGND _06154_ sg13g2_a21oi_1
X_25887_ _04338_ _06151_ _06154_ VPWR VGND _06155_ sg13g2_a21oi_1
X_25888_ _00120_ _03733_ _03737_ _02437_ _06155_ VPWR 
+ VGND
+ _06156_ sg13g2_a221oi_1
X_25889_ _04357_ _02138_ VPWR VGND _06157_ sg13g2_nor2_1
X_25890_ _02161_ _03881_ VPWR VGND _06158_ sg13g2_nor2_1
X_25891_ _04662_ _06157_ _06158_ _04362_ VPWR VGND 
+ _06159_
+ sg13g2_a22oi_1
X_25892_ _02138_ _03907_ VPWR VGND _06160_ sg13g2_nand2b_1
X_25893_ _04365_ _02161_ _06160_ VPWR VGND _06161_ sg13g2_o21ai_1
X_25894_ _04666_ _06161_ _04021_ VPWR VGND _06162_ sg13g2_a21oi_1
X_25895_ _04355_ _06159_ _06162_ VPWR VGND _06163_ sg13g2_a21oi_1
X_25896_ _00121_ _04353_ _04354_ _02188_ _06163_ VPWR 
+ VGND
+ _06164_ sg13g2_a221oi_1
X_25897_ _04337_ _06156_ _06164_ _04330_ _04688_ VPWR 
+ VGND
+ _06165_ sg13g2_a221oi_1
X_25898_ _02713_ _02621_ VPWR VGND _06166_ sg13g2_nor2_1
X_25899_ _02642_ _04533_ VPWR VGND _06167_ sg13g2_nor2_1
X_25900_ _04568_ _06166_ _06167_ _04536_ VPWR VGND 
+ _06168_
+ sg13g2_a22oi_1
X_25901_ _02621_ _04320_ VPWR VGND _06169_ sg13g2_nand2b_1
X_25902_ _03887_ _02642_ _06169_ VPWR VGND _06170_ sg13g2_o21ai_1
X_25903_ _04573_ _06170_ _04542_ VPWR VGND _06171_ sg13g2_a21oi_1
X_25904_ _04530_ _06168_ _06171_ VPWR VGND _06172_ sg13g2_a21oi_1
X_25905_ _00119_ _04660_ _04661_ _02667_ _06172_ VPWR 
+ VGND
+ _06173_ sg13g2_a221oi_1
X_25906_ _05483_ _06173_ VPWR VGND _06174_ sg13g2_nand2_1
X_25907_ \atbs_core_0.spike_memory_0.n2385_o[3]\ _03735_ VPWR VGND _06175_ sg13g2_nand2b_1
X_25908_ \atbs_core_0.spike_memory_0.n2382_o[3]\ _04102_ _06175_ VPWR VGND _06176_ sg13g2_o21ai_1
X_25909_ _04346_ _02289_ VPWR VGND _06177_ sg13g2_nor2_1
X_25910_ _02313_ _04265_ VPWR VGND _06178_ sg13g2_nor2_1
X_25911_ _05496_ _06177_ _06178_ _04112_ VPWR VGND 
+ _06179_
+ sg13g2_a22oi_1
X_25912_ _02289_ _03760_ VPWR VGND _06180_ sg13g2_nand2b_1
X_25913_ _04267_ _02313_ _06180_ VPWR VGND _06181_ sg13g2_o21ai_1
X_25914_ _04235_ _06181_ _03973_ VPWR VGND _06182_ sg13g2_a21oi_1
X_25915_ _03940_ _06179_ _06182_ VPWR VGND _06183_ sg13g2_a21oi_1
X_25916_ _06176_ _06183_ VPWR VGND _06184_ sg13g2_or2_1
X_25917_ \atbs_core_0.spike_memory_0.n2381_o[3]\ _04075_ VPWR VGND _06185_ sg13g2_nor2_1
X_25918_ \atbs_core_0.spike_memory_0.n2378_o[3]\ _04229_ VPWR VGND _06186_ sg13g2_nor2_1
X_25919_ _04480_ _02235_ VPWR VGND _06187_ sg13g2_nor2_1
X_25920_ _02258_ _03742_ VPWR VGND _06188_ sg13g2_nor2_1
X_25921_ _04422_ _06187_ _06188_ _03827_ VPWR VGND 
+ _06189_
+ sg13g2_a22oi_1
X_25922_ _02235_ _04050_ VPWR VGND _06190_ sg13g2_nand2b_1
X_25923_ _03915_ _02258_ _06190_ VPWR VGND _06191_ sg13g2_o21ai_1
X_25924_ _05510_ _06191_ _03738_ VPWR VGND _06192_ sg13g2_a21oi_1
X_25925_ _04839_ _06189_ _06192_ VPWR VGND _06193_ sg13g2_a21oi_1
X_25926_ _03773_ _06185_ _06186_ _06193_ VPWR VGND 
+ _06194_
+ sg13g2_nor4_1
X_25927_ \atbs_core_0.spike_memory_0.n2389_o[3]\ _04759_ VPWR VGND _06195_ sg13g2_nor2_1
X_25928_ \atbs_core_0.spike_memory_0.n2386_o[3]\ _04000_ VPWR VGND _06196_ sg13g2_nor2_1
X_25929_ _03863_ _02345_ VPWR VGND _06197_ sg13g2_nor2_1
X_25930_ _02369_ _05245_ VPWR VGND _06198_ sg13g2_nor2_1
X_25931_ _04086_ _06197_ _06198_ _03864_ VPWR VGND 
+ _06199_
+ sg13g2_a22oi_1
X_25932_ _02345_ _03854_ VPWR VGND _06200_ sg13g2_nand2b_1
X_25933_ _04480_ _02369_ _06200_ VPWR VGND _06201_ sg13g2_o21ai_1
X_25934_ _05510_ _06201_ _03810_ VPWR VGND _06202_ sg13g2_a21oi_1
X_25935_ _04098_ _06199_ _06202_ VPWR VGND _06203_ sg13g2_a21oi_1
X_25936_ _04746_ _06195_ _06196_ _06203_ VPWR VGND 
+ _06204_
+ sg13g2_nor4_1
X_25937_ _06194_ _06204_ _03924_ VPWR VGND _06205_ sg13g2_o21ai_1
X_25938_ _04277_ _06184_ _06205_ VPWR VGND _06206_ sg13g2_o21ai_1
X_25939_ \atbs_core_0.spike_memory_0.n2405_o[3]\ _04245_ VPWR VGND _06207_ sg13g2_nor2_1
X_25940_ \atbs_core_0.spike_memory_0.n2402_o[3]\ _04247_ VPWR VGND _06208_ sg13g2_nor2_1
X_25941_ _04413_ _02574_ VPWR VGND _06209_ sg13g2_nor2_1
X_25942_ _02595_ _04422_ VPWR VGND _06210_ sg13g2_nor2_1
X_25943_ _04280_ _06209_ _06210_ _04704_ VPWR VGND 
+ _06211_
+ sg13g2_a22oi_1
X_25944_ _02574_ _04425_ VPWR VGND _06212_ sg13g2_nand2b_1
X_25945_ _05533_ _02595_ _06212_ VPWR VGND _06213_ sg13g2_o21ai_1
X_25946_ _04092_ _06213_ _04839_ VPWR VGND _06214_ sg13g2_a21oi_1
X_25947_ _03769_ _06211_ _06214_ VPWR VGND _06215_ sg13g2_a21oi_1
X_25948_ _12094_ _06207_ _06208_ _06215_ VPWR VGND 
+ _06216_
+ sg13g2_nor4_1
X_25949_ \atbs_core_0.spike_memory_0.n2401_o[3]\ _04372_ VPWR VGND _06217_ sg13g2_nor2_1
X_25950_ \atbs_core_0.spike_memory_0.n2398_o[3]\ _05540_ _03723_ VPWR VGND _06218_ sg13g2_o21ai_1
X_25951_ _04026_ _02526_ VPWR VGND _06219_ sg13g2_nor2_1
X_25952_ _02548_ _03975_ VPWR VGND _06220_ sg13g2_nor2_1
X_25953_ _04152_ _06219_ _06220_ _05544_ VPWR VGND 
+ _06221_
+ sg13g2_a22oi_1
X_25954_ _02526_ _04115_ VPWR VGND _06222_ sg13g2_nand2b_1
X_25955_ _03764_ _02548_ _06222_ VPWR VGND _06223_ sg13g2_o21ai_1
X_25956_ _04114_ _06223_ _04118_ VPWR VGND _06224_ sg13g2_a21oi_1
X_25957_ _04142_ _06221_ _06224_ VPWR VGND _06225_ sg13g2_a21oi_1
X_25958_ _06217_ _06218_ _06225_ VPWR VGND _06226_ sg13g2_nor3_1
X_25959_ \atbs_core_0.spike_memory_0.n2397_o[3]\ _04260_ VPWR VGND _06227_ sg13g2_nor2_1
X_25960_ \atbs_core_0.spike_memory_0.n2394_o[3]\ _04079_ VPWR VGND _06228_ sg13g2_nor2_1
X_25961_ _04236_ _02478_ VPWR VGND _06229_ sg13g2_nor2_1
X_25962_ _02500_ _04250_ VPWR VGND _06230_ sg13g2_nor2_1
X_25963_ _03884_ _06229_ _06230_ _04268_ VPWR VGND 
+ _06231_
+ sg13g2_a22oi_1
X_25964_ _02478_ _04004_ VPWR VGND _06232_ sg13g2_nand2b_1
X_25965_ _04083_ _02500_ _06232_ VPWR VGND _06233_ sg13g2_o21ai_1
X_25966_ _04253_ _06233_ _04272_ VPWR VGND _06234_ sg13g2_a21oi_1
X_25967_ _04263_ _06231_ _06234_ VPWR VGND _06235_ sg13g2_a21oi_1
X_25968_ _04244_ _06227_ _06228_ _06235_ VPWR VGND 
+ _06236_
+ sg13g2_nor4_1
X_25969_ _06216_ _06226_ _06236_ VPWR VGND _06237_ sg13g2_or3_1
X_25970_ _04330_ _06206_ _06237_ _03718_ _04336_ VPWR 
+ VGND
+ _06238_ sg13g2_a221oi_1
X_25971_ \atbs_core_0.spike_memory_0.n2413_o[3]\ _04372_ VPWR VGND _06239_ sg13g2_nor2_1
X_25972_ \atbs_core_0.spike_memory_0.n2410_o[3]\ _04527_ VPWR VGND _06240_ sg13g2_nor2_1
X_25973_ _03747_ _12520_ VPWR VGND _06241_ sg13g2_nor2_1
X_25974_ _12543_ _03751_ VPWR VGND _06242_ sg13g2_nor2_1
X_25975_ _03744_ _06241_ _06242_ _04379_ VPWR VGND 
+ _06243_
+ sg13g2_a22oi_1
X_25976_ _12520_ _03764_ VPWR VGND _06244_ sg13g2_nand2b_1
X_25977_ _04512_ _12543_ _06244_ VPWR VGND _06245_ sg13g2_o21ai_1
X_25978_ _04387_ _06245_ _04392_ VPWR VGND _06246_ sg13g2_a21oi_1
X_25979_ _03740_ _06243_ _06246_ VPWR VGND _06247_ sg13g2_a21oi_1
X_25980_ _03800_ _06239_ _06240_ _06247_ VPWR VGND 
+ _06248_
+ sg13g2_nor4_1
X_25981_ \atbs_core_0.spike_memory_0.n2417_o[3]\ _03944_ VPWR VGND _06249_ sg13g2_nor2_1
X_25982_ \atbs_core_0.spike_memory_0.n2414_o[3]\ _04032_ _03966_ VPWR VGND _06250_ sg13g2_o21ai_1
X_25983_ _03822_ _12575_ VPWR VGND _06251_ sg13g2_nor2_1
X_25984_ _12599_ _03909_ VPWR VGND _06252_ sg13g2_nor2_1
X_25985_ _03906_ _06251_ _06252_ _03911_ VPWR VGND 
+ _06253_
+ sg13g2_a22oi_1
X_25986_ _12575_ _05745_ VPWR VGND _06254_ sg13g2_nand2b_1
X_25987_ _03914_ _12599_ _06254_ VPWR VGND _06255_ sg13g2_o21ai_1
X_25988_ _03913_ _06255_ _03919_ VPWR VGND _06256_ sg13g2_a21oi_1
X_25989_ _03905_ _06253_ _06256_ VPWR VGND _06257_ sg13g2_a21oi_1
X_25990_ _06249_ _06250_ _06257_ VPWR VGND _06258_ sg13g2_nor3_1
X_25991_ \atbs_core_0.spike_memory_0.n2436_q[1200]\ _03877_ VPWR VGND _06259_ sg13g2_nor2_1
X_25992_ \atbs_core_0.spike_memory_0.n2418_o[3]\ _04702_ VPWR VGND _06260_ sg13g2_nor2_1
X_25993_ _05753_ _12633_ VPWR VGND _06261_ sg13g2_nor2_1
X_25994_ _12658_ _05496_ VPWR VGND _06262_ sg13g2_nor2_1
X_25995_ _04628_ _06261_ _06262_ _02713_ VPWR VGND 
+ _06263_
+ sg13g2_a22oi_1
X_25996_ _12633_ _03892_ VPWR VGND _06264_ sg13g2_nand2b_1
X_25997_ _02712_ _12658_ _06264_ VPWR VGND _06265_ sg13g2_o21ai_1
X_25998_ _03889_ _06265_ _04263_ VPWR VGND _06266_ sg13g2_a21oi_1
X_25999_ _04635_ _06263_ _06266_ VPWR VGND _06267_ sg13g2_a21oi_1
X_26000_ _12095_ _06259_ _06260_ _06267_ VPWR VGND 
+ _06268_
+ sg13g2_nor4_1
X_26001_ _06248_ _06258_ _06268_ VPWR VGND _06269_ sg13g2_nor3_1
X_26002_ _06269_ _05483_ VPWR VGND _06270_ sg13g2_nand2b_1
X_26003_ _06165_ _06174_ _06238_ _06270_ VPWR VGND 
+ _06271_
+ sg13g2_a22oi_1
X_26004_ \atbs_core_0.spike_memory_0.n2361_o[3]\ _04373_ VPWR VGND _06272_ sg13g2_nor2_1
X_26005_ \atbs_core_0.spike_memory_0.n2358_o[3]\ _04508_ VPWR VGND _06273_ sg13g2_nor2_1
X_26006_ _04513_ _02073_ VPWR VGND _06274_ sg13g2_nor2_1
X_26007_ _02256_ _04716_ VPWR VGND _06275_ sg13g2_nor2_1
X_26008_ _04511_ _06274_ _06275_ _04613_ VPWR VGND 
+ _06276_
+ sg13g2_a22oi_1
X_26009_ _02073_ _04518_ VPWR VGND _06277_ sg13g2_nand2b_1
X_26010_ _04383_ _02256_ _06277_ VPWR VGND _06278_ sg13g2_o21ai_1
X_26011_ _04517_ _06278_ _04521_ VPWR VGND _06279_ sg13g2_a21oi_1
X_26012_ _04608_ _06276_ _06279_ VPWR VGND _06280_ sg13g2_a21oi_1
X_26013_ _04505_ _06272_ _06273_ _06280_ VPWR VGND 
+ _06281_
+ sg13g2_nor4_1
X_26014_ \atbs_core_0.spike_memory_0.n2369_o[3]\ _04525_ VPWR VGND _06282_ sg13g2_nor2_1
X_26015_ \atbs_core_0.spike_memory_0.n2366_o[3]\ _04549_ VPWR VGND _06283_ sg13g2_nor2_1
X_26016_ _04553_ _02029_ VPWR VGND _06284_ sg13g2_nor2_1
X_26017_ _02050_ _04533_ VPWR VGND _06285_ sg13g2_nor2_1
X_26018_ _04531_ _06284_ _06285_ _04557_ VPWR VGND 
+ _06286_
+ sg13g2_a22oi_1
X_26019_ _02029_ _04559_ VPWR VGND _06287_ sg13g2_nand2b_1
X_26020_ _04539_ _02050_ _06287_ VPWR VGND _06288_ sg13g2_o21ai_1
X_26021_ _04538_ _06288_ _04562_ VPWR VGND _06289_ sg13g2_a21oi_1
X_26022_ _04551_ _06286_ _06289_ VPWR VGND _06290_ sg13g2_a21oi_1
X_26023_ _04604_ _06282_ _06283_ _06290_ VPWR VGND 
+ _06291_
+ sg13g2_nor4_1
X_26024_ _04504_ _06281_ _06291_ VPWR VGND _06292_ sg13g2_nor3_1
X_26025_ \atbs_core_0.spike_memory_0.n2365_o[3]\ _04506_ VPWR VGND _06293_ sg13g2_nor2_1
X_26026_ \atbs_core_0.spike_memory_0.n2362_o[3]\ _04508_ VPWR VGND _06294_ sg13g2_nor2_1
X_26027_ _04535_ _12656_ VPWR VGND _06295_ sg13g2_nor2_1
X_26028_ _12655_ _04555_ VPWR VGND _06296_ sg13g2_nor2_1
X_26029_ _04378_ _06295_ _06296_ _04557_ VPWR VGND 
+ _06297_
+ sg13g2_a22oi_1
X_26030_ _12656_ _05544_ VPWR VGND _06298_ sg13g2_nand2b_1
X_26031_ _03755_ _12655_ _06298_ VPWR VGND _06299_ sg13g2_o21ai_1
X_26032_ _04388_ _06299_ _04562_ VPWR VGND _06300_ sg13g2_a21oi_1
X_26033_ _04551_ _06297_ _06300_ VPWR VGND _06301_ sg13g2_a21oi_1
X_26034_ _03968_ _06293_ _06294_ _06301_ VPWR VGND 
+ _06302_
+ sg13g2_nor4_1
X_26035_ \atbs_core_0.spike_memory_0.n2373_o[3]\ _12088_ VPWR VGND _06303_ sg13g2_nor2_1
X_26036_ \atbs_core_0.spike_memory_0.n2370_o[3]\ _04528_ VPWR VGND _06304_ sg13g2_nor2_1
X_26037_ _03934_ _02083_ VPWR VGND _06305_ sg13g2_nor2_1
X_26038_ _02105_ _04570_ VPWR VGND _06306_ sg13g2_nor2_1
X_26039_ _04568_ _06305_ _06306_ _02714_ VPWR VGND 
+ _06307_
+ sg13g2_a22oi_1
X_26040_ _02083_ _04361_ VPWR VGND _06308_ sg13g2_nand2b_1
X_26041_ _04574_ _02105_ _06308_ VPWR VGND _06309_ sg13g2_o21ai_1
X_26042_ _04573_ _06309_ _04338_ VPWR VGND _06310_ sg13g2_a21oi_1
X_26043_ _02702_ _06307_ _06310_ VPWR VGND _06311_ sg13g2_a21oi_1
X_26044_ _04126_ _06303_ _06304_ _06311_ VPWR VGND 
+ _06312_
+ sg13g2_nor4_1
X_26045_ _04547_ _06302_ _06312_ VPWR VGND _06313_ sg13g2_nor3_1
X_26046_ _07549_ _06292_ _06313_ VPWR VGND _06314_ sg13g2_nor3_1
X_26047_ _04333_ _06271_ _06314_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[3]\ sg13g2_a21o_1
X_26048_ _04340_ _02396_ VPWR VGND _06315_ sg13g2_nor2_1
X_26049_ _02415_ _03976_ VPWR VGND _06316_ sg13g2_nor2_1
X_26050_ _04339_ _06315_ _06316_ _04343_ VPWR VGND 
+ _06317_
+ sg13g2_a22oi_1
X_26051_ _02396_ _03788_ VPWR VGND _06318_ sg13g2_nand2b_1
X_26052_ _04347_ _02415_ _06318_ VPWR VGND _06319_ sg13g2_o21ai_1
X_26053_ _04345_ _06319_ _04684_ VPWR VGND _06320_ sg13g2_a21oi_1
X_26054_ _04338_ _06317_ _06320_ VPWR VGND _06321_ sg13g2_a21oi_1
X_26055_ _00123_ _03733_ _03737_ _02439_ _06321_ VPWR 
+ VGND
+ _06322_ sg13g2_a221oi_1
X_26056_ _04357_ _02139_ VPWR VGND _06323_ sg13g2_nor2_1
X_26057_ _02162_ _04359_ VPWR VGND _06324_ sg13g2_nor2_1
X_26058_ _04356_ _06323_ _06324_ _04362_ VPWR VGND 
+ _06325_
+ sg13g2_a22oi_1
X_26059_ _02139_ _03907_ VPWR VGND _06326_ sg13g2_nand2b_1
X_26060_ _04365_ _02162_ _06326_ VPWR VGND _06327_ sg13g2_o21ai_1
X_26061_ _04364_ _06327_ _04021_ VPWR VGND _06328_ sg13g2_a21oi_1
X_26062_ _04355_ _06325_ _06328_ VPWR VGND _06329_ sg13g2_a21oi_1
X_26063_ _00124_ _04353_ _04354_ _02190_ _06329_ VPWR 
+ VGND
+ _06330_ sg13g2_a221oi_1
X_26064_ _04337_ _06322_ _06330_ _04371_ _04688_ VPWR 
+ VGND
+ _06331_ sg13g2_a221oi_1
X_26065_ _02713_ _02622_ VPWR VGND _06332_ sg13g2_nor2_1
X_26066_ _02643_ _04533_ VPWR VGND _06333_ sg13g2_nor2_1
X_26067_ _04531_ _06332_ _06333_ _04536_ VPWR VGND 
+ _06334_
+ sg13g2_a22oi_1
X_26068_ _02622_ _04320_ VPWR VGND _06335_ sg13g2_nand2b_1
X_26069_ _03887_ _02643_ _06335_ VPWR VGND _06336_ sg13g2_o21ai_1
X_26070_ _04538_ _06336_ _04542_ VPWR VGND _06337_ sg13g2_a21oi_1
X_26071_ _04530_ _06334_ _06337_ VPWR VGND _06338_ sg13g2_a21oi_1
X_26072_ _00122_ _04660_ _04661_ _02669_ _06338_ VPWR 
+ VGND
+ _06339_ sg13g2_a221oi_1
X_26073_ _05483_ _06339_ VPWR VGND _06340_ sg13g2_nand2_1
X_26074_ \atbs_core_0.spike_memory_0.n2385_o[4]\ _03735_ VPWR VGND _06341_ sg13g2_nand2b_1
X_26075_ \atbs_core_0.spike_memory_0.n2382_o[4]\ _04102_ _06341_ VPWR VGND _06342_ sg13g2_o21ai_1
X_26076_ _04346_ _02291_ VPWR VGND _06343_ sg13g2_nor2_1
X_26077_ _02314_ _04265_ VPWR VGND _06344_ sg13g2_nor2_1
X_26078_ _05496_ _06343_ _06344_ _04112_ VPWR VGND 
+ _06345_
+ sg13g2_a22oi_1
X_26079_ _02291_ _03760_ VPWR VGND _06346_ sg13g2_nand2b_1
X_26080_ _04267_ _02314_ _06346_ VPWR VGND _06347_ sg13g2_o21ai_1
X_26081_ _04235_ _06347_ _03973_ VPWR VGND _06348_ sg13g2_a21oi_1
X_26082_ _03940_ _06345_ _06348_ VPWR VGND _06349_ sg13g2_a21oi_1
X_26083_ _06342_ _06349_ VPWR VGND _06350_ sg13g2_or2_1
X_26084_ \atbs_core_0.spike_memory_0.n2381_o[4]\ _04075_ VPWR VGND _06351_ sg13g2_nor2_1
X_26085_ \atbs_core_0.spike_memory_0.n2378_o[4]\ _04229_ VPWR VGND _06352_ sg13g2_nor2_1
X_26086_ _04480_ _02236_ VPWR VGND _06353_ sg13g2_nor2_1
X_26087_ _02259_ _03742_ VPWR VGND _06354_ sg13g2_nor2_1
X_26088_ _04422_ _06353_ _06354_ _03827_ VPWR VGND 
+ _06355_
+ sg13g2_a22oi_1
X_26089_ _02236_ _03745_ VPWR VGND _06356_ sg13g2_nand2b_1
X_26090_ _03915_ _02259_ _06356_ VPWR VGND _06357_ sg13g2_o21ai_1
X_26091_ _05510_ _06357_ _03738_ VPWR VGND _06358_ sg13g2_a21oi_1
X_26092_ _04839_ _06355_ _06358_ VPWR VGND _06359_ sg13g2_a21oi_1
X_26093_ _03773_ _06351_ _06352_ _06359_ VPWR VGND 
+ _06360_
+ sg13g2_nor4_1
X_26094_ \atbs_core_0.spike_memory_0.n2389_o[4]\ _04075_ VPWR VGND _06361_ sg13g2_nor2_1
X_26095_ \atbs_core_0.spike_memory_0.n2386_o[4]\ _04000_ VPWR VGND _06362_ sg13g2_nor2_1
X_26096_ _03863_ _02346_ VPWR VGND _06363_ sg13g2_nor2_1
X_26097_ _02370_ _05245_ VPWR VGND _06364_ sg13g2_nor2_1
X_26098_ _04086_ _06363_ _06364_ _04167_ VPWR VGND 
+ _06365_
+ sg13g2_a22oi_1
X_26099_ _02346_ _03854_ VPWR VGND _06366_ sg13g2_nand2b_1
X_26100_ _04480_ _02370_ _06366_ VPWR VGND _06367_ sg13g2_o21ai_1
X_26101_ _05510_ _06367_ _03738_ VPWR VGND _06368_ sg13g2_a21oi_1
X_26102_ _04098_ _06365_ _06368_ VPWR VGND _06369_ sg13g2_a21oi_1
X_26103_ _04746_ _06361_ _06362_ _06369_ VPWR VGND 
+ _06370_
+ sg13g2_nor4_1
X_26104_ _06360_ _06370_ _03924_ VPWR VGND _06371_ sg13g2_o21ai_1
X_26105_ _04277_ _06350_ _06371_ VPWR VGND _06372_ sg13g2_o21ai_1
X_26106_ \atbs_core_0.spike_memory_0.n2405_o[4]\ _04245_ VPWR VGND _06373_ sg13g2_nor2_1
X_26107_ \atbs_core_0.spike_memory_0.n2402_o[4]\ _04247_ VPWR VGND _06374_ sg13g2_nor2_1
X_26108_ _04413_ _02575_ VPWR VGND _06375_ sg13g2_nor2_1
X_26109_ _02596_ _04422_ VPWR VGND _06376_ sg13g2_nor2_1
X_26110_ _04280_ _06375_ _06376_ _04704_ VPWR VGND 
+ _06377_
+ sg13g2_a22oi_1
X_26111_ _02575_ _04425_ VPWR VGND _06378_ sg13g2_nand2b_1
X_26112_ _05533_ _02596_ _06378_ VPWR VGND _06379_ sg13g2_o21ai_1
X_26113_ _04092_ _06379_ _04287_ VPWR VGND _06380_ sg13g2_a21oi_1
X_26114_ _03769_ _06377_ _06380_ VPWR VGND _06381_ sg13g2_a21oi_1
X_26115_ _12094_ _06373_ _06374_ _06381_ VPWR VGND 
+ _06382_
+ sg13g2_nor4_1
X_26116_ \atbs_core_0.spike_memory_0.n2401_o[4]\ _04076_ VPWR VGND _06383_ sg13g2_nor2_1
X_26117_ \atbs_core_0.spike_memory_0.n2398_o[4]\ _05540_ _03723_ VPWR VGND _06384_ sg13g2_o21ai_1
X_26118_ _04026_ _02527_ VPWR VGND _06385_ sg13g2_nor2_1
X_26119_ _02549_ _03975_ VPWR VGND _06386_ sg13g2_nor2_1
X_26120_ _04152_ _06385_ _06386_ _05544_ VPWR VGND 
+ _06387_
+ sg13g2_a22oi_1
X_26121_ _02527_ _04115_ VPWR VGND _06388_ sg13g2_nand2b_1
X_26122_ _03764_ _02549_ _06388_ VPWR VGND _06389_ sg13g2_o21ai_1
X_26123_ _04114_ _06389_ _04118_ VPWR VGND _06390_ sg13g2_a21oi_1
X_26124_ _04142_ _06387_ _06390_ VPWR VGND _06391_ sg13g2_a21oi_1
X_26125_ _06383_ _06384_ _06391_ VPWR VGND _06392_ sg13g2_nor3_1
X_26126_ \atbs_core_0.spike_memory_0.n2397_o[4]\ _04260_ VPWR VGND _06393_ sg13g2_nor2_1
X_26127_ \atbs_core_0.spike_memory_0.n2394_o[4]\ _04079_ VPWR VGND _06394_ sg13g2_nor2_1
X_26128_ _04236_ _02479_ VPWR VGND _06395_ sg13g2_nor2_1
X_26129_ _02501_ _04250_ VPWR VGND _06396_ sg13g2_nor2_1
X_26130_ _03884_ _06395_ _06396_ _04268_ VPWR VGND 
+ _06397_
+ sg13g2_a22oi_1
X_26131_ _02479_ _04004_ VPWR VGND _06398_ sg13g2_nand2b_1
X_26132_ _04083_ _02501_ _06398_ VPWR VGND _06399_ sg13g2_o21ai_1
X_26133_ _04253_ _06399_ _04272_ VPWR VGND _06400_ sg13g2_a21oi_1
X_26134_ _03895_ _06397_ _06400_ VPWR VGND _06401_ sg13g2_a21oi_1
X_26135_ _04244_ _06393_ _06394_ _06401_ VPWR VGND 
+ _06402_
+ sg13g2_nor4_1
X_26136_ _06382_ _06392_ _06402_ VPWR VGND _06403_ sg13g2_or3_1
X_26137_ _04330_ _06372_ _06403_ _03718_ _04336_ VPWR 
+ VGND
+ _06404_ sg13g2_a221oi_1
X_26138_ \atbs_core_0.spike_memory_0.n2413_o[4]\ _04372_ VPWR VGND _06405_ sg13g2_nor2_1
X_26139_ \atbs_core_0.spike_memory_0.n2410_o[4]\ _04527_ VPWR VGND _06406_ sg13g2_nor2_1
X_26140_ _03747_ _12521_ VPWR VGND _06407_ sg13g2_nor2_1
X_26141_ _12545_ _03751_ VPWR VGND _06408_ sg13g2_nor2_1
X_26142_ _03744_ _06407_ _06408_ _04379_ VPWR VGND 
+ _06409_
+ sg13g2_a22oi_1
X_26143_ _12521_ _04111_ VPWR VGND _06410_ sg13g2_nand2b_1
X_26144_ _04512_ _12545_ _06410_ VPWR VGND _06411_ sg13g2_o21ai_1
X_26145_ _04387_ _06411_ _04392_ VPWR VGND _06412_ sg13g2_a21oi_1
X_26146_ _04376_ _06409_ _06412_ VPWR VGND _06413_ sg13g2_a21oi_1
X_26147_ _03800_ _06405_ _06406_ _06413_ VPWR VGND 
+ _06414_
+ sg13g2_nor4_1
X_26148_ \atbs_core_0.spike_memory_0.n2417_o[4]\ _03944_ VPWR VGND _06415_ sg13g2_nor2_1
X_26149_ \atbs_core_0.spike_memory_0.n2414_o[4]\ _04230_ _03723_ VPWR VGND _06416_ sg13g2_o21ai_1
X_26150_ _03822_ _12576_ VPWR VGND _06417_ sg13g2_nor2_1
X_26151_ _12600_ _03909_ VPWR VGND _06418_ sg13g2_nor2_1
X_26152_ _03906_ _06417_ _06418_ _03911_ VPWR VGND 
+ _06419_
+ sg13g2_a22oi_1
X_26153_ _12576_ _05745_ VPWR VGND _06420_ sg13g2_nand2b_1
X_26154_ _03914_ _12600_ _06420_ VPWR VGND _06421_ sg13g2_o21ai_1
X_26155_ _03913_ _06421_ _03919_ VPWR VGND _06422_ sg13g2_a21oi_1
X_26156_ _03905_ _06419_ _06422_ VPWR VGND _06423_ sg13g2_a21oi_1
X_26157_ _06415_ _06416_ _06423_ VPWR VGND _06424_ sg13g2_nor3_1
X_26158_ \atbs_core_0.spike_memory_0.n2436_q[1201]\ _03877_ VPWR VGND _06425_ sg13g2_nor2_1
X_26159_ \atbs_core_0.spike_memory_0.n2418_o[4]\ _04702_ VPWR VGND _06426_ sg13g2_nor2_1
X_26160_ _05753_ _12634_ VPWR VGND _06427_ sg13g2_nor2_1
X_26161_ _12659_ _05496_ VPWR VGND _06428_ sg13g2_nor2_1
X_26162_ _04628_ _06427_ _06428_ _02713_ VPWR VGND 
+ _06429_
+ sg13g2_a22oi_1
X_26163_ _12634_ _03892_ VPWR VGND _06430_ sg13g2_nand2b_1
X_26164_ _03882_ _12659_ _06430_ VPWR VGND _06431_ sg13g2_o21ai_1
X_26165_ _03889_ _06431_ _04263_ VPWR VGND _06432_ sg13g2_a21oi_1
X_26166_ _04635_ _06429_ _06432_ VPWR VGND _06433_ sg13g2_a21oi_1
X_26167_ _12095_ _06425_ _06426_ _06433_ VPWR VGND 
+ _06434_
+ sg13g2_nor4_1
X_26168_ _06414_ _06424_ _06434_ VPWR VGND _06435_ sg13g2_nor3_1
X_26169_ _06435_ _05483_ VPWR VGND _06436_ sg13g2_nand2b_1
X_26170_ _06331_ _06340_ _06404_ _06436_ VPWR VGND 
+ _06437_
+ sg13g2_a22oi_1
X_26171_ \atbs_core_0.spike_memory_0.n2361_o[4]\ _04373_ VPWR VGND _06438_ sg13g2_nor2_1
X_26172_ \atbs_core_0.spike_memory_0.n2358_o[4]\ _04508_ VPWR VGND _06439_ sg13g2_nor2_1
X_26173_ _04513_ _02077_ VPWR VGND _06440_ sg13g2_nor2_1
X_26174_ _02268_ _04716_ VPWR VGND _06441_ sg13g2_nor2_1
X_26175_ _04511_ _06440_ _06441_ _04613_ VPWR VGND 
+ _06442_
+ sg13g2_a22oi_1
X_26176_ _02077_ _04518_ VPWR VGND _06443_ sg13g2_nand2b_1
X_26177_ _03984_ _02268_ _06443_ VPWR VGND _06444_ sg13g2_o21ai_1
X_26178_ _04517_ _06444_ _04521_ VPWR VGND _06445_ sg13g2_a21oi_1
X_26179_ _04608_ _06442_ _06445_ VPWR VGND _06446_ sg13g2_a21oi_1
X_26180_ _04505_ _06438_ _06439_ _06446_ VPWR VGND 
+ _06447_
+ sg13g2_nor4_1
X_26181_ \atbs_core_0.spike_memory_0.n2369_o[4]\ _04525_ VPWR VGND _06448_ sg13g2_nor2_1
X_26182_ \atbs_core_0.spike_memory_0.n2366_o[4]\ _04549_ VPWR VGND _06449_ sg13g2_nor2_1
X_26183_ _04553_ _02030_ VPWR VGND _06450_ sg13g2_nor2_1
X_26184_ _02051_ _04533_ VPWR VGND _06451_ sg13g2_nor2_1
X_26185_ _04531_ _06450_ _06451_ _04557_ VPWR VGND 
+ _06452_
+ sg13g2_a22oi_1
X_26186_ _02030_ _04559_ VPWR VGND _06453_ sg13g2_nand2b_1
X_26187_ _04539_ _02051_ _06453_ VPWR VGND _06454_ sg13g2_o21ai_1
X_26188_ _04538_ _06454_ _04562_ VPWR VGND _06455_ sg13g2_a21oi_1
X_26189_ _04551_ _06452_ _06455_ VPWR VGND _06456_ sg13g2_a21oi_1
X_26190_ _04604_ _06448_ _06449_ _06456_ VPWR VGND 
+ _06457_
+ sg13g2_nor4_1
X_26191_ _03925_ _06447_ _06457_ VPWR VGND _06458_ sg13g2_nor3_1
X_26192_ \atbs_core_0.spike_memory_0.n2365_o[4]\ _04506_ VPWR VGND _06459_ sg13g2_nor2_1
X_26193_ \atbs_core_0.spike_memory_0.n2362_o[4]\ _04508_ VPWR VGND _06460_ sg13g2_nor2_1
X_26194_ _04535_ _12669_ VPWR VGND _06461_ sg13g2_nor2_1
X_26195_ _12668_ _04555_ VPWR VGND _06462_ sg13g2_nor2_1
X_26196_ _04378_ _06461_ _06462_ _04557_ VPWR VGND 
+ _06463_
+ sg13g2_a22oi_1
X_26197_ _12669_ _05544_ VPWR VGND _06464_ sg13g2_nand2b_1
X_26198_ _03755_ _12668_ _06464_ VPWR VGND _06465_ sg13g2_o21ai_1
X_26199_ _04388_ _06465_ _04393_ VPWR VGND _06466_ sg13g2_a21oi_1
X_26200_ _04551_ _06463_ _06466_ VPWR VGND _06467_ sg13g2_a21oi_1
X_26201_ _03968_ _06459_ _06460_ _06467_ VPWR VGND 
+ _06468_
+ sg13g2_nor4_1
X_26202_ \atbs_core_0.spike_memory_0.n2373_o[4]\ _12088_ VPWR VGND _06469_ sg13g2_nor2_1
X_26203_ \atbs_core_0.spike_memory_0.n2370_o[4]\ _04528_ VPWR VGND _06470_ sg13g2_nor2_1
X_26204_ _03934_ _02084_ VPWR VGND _06471_ sg13g2_nor2_1
X_26205_ _02107_ _04570_ VPWR VGND _06472_ sg13g2_nor2_1
X_26206_ _04568_ _06471_ _06472_ _02714_ VPWR VGND 
+ _06473_
+ sg13g2_a22oi_1
X_26207_ _02084_ _04361_ VPWR VGND _06474_ sg13g2_nand2b_1
X_26208_ _04574_ _02107_ _06474_ VPWR VGND _06475_ sg13g2_o21ai_1
X_26209_ _04573_ _06475_ _04542_ VPWR VGND _06476_ sg13g2_a21oi_1
X_26210_ _02702_ _06473_ _06476_ VPWR VGND _06477_ sg13g2_a21oi_1
X_26211_ _04126_ _06469_ _06470_ _06477_ VPWR VGND 
+ _06478_
+ sg13g2_nor4_1
X_26212_ _04547_ _06468_ _06478_ VPWR VGND _06479_ sg13g2_nor3_1
X_26213_ _07549_ _06458_ _06479_ VPWR VGND _06480_ sg13g2_nor3_1
X_26214_ _04503_ _06437_ _06480_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[4]\ sg13g2_a21o_1
X_26215_ \atbs_core_0.spike_memory_0.n2392_o[5]\ _04387_ VPWR VGND _06481_ sg13g2_nand2_1
X_26216_ _00126_ _03861_ _06481_ VPWR VGND _06482_ sg13g2_o21ai_1
X_26217_ \atbs_core_0.spike_memory_0.n2391_o[5]\ _06068_ _06482_ _07561_ VPWR VGND 
+ _06483_
+ sg13g2_a22oi_1
X_26218_ _02441_ _12088_ _06483_ VPWR VGND _06484_ sg13g2_o21ai_1
X_26219_ _04357_ _02140_ VPWR VGND _06485_ sg13g2_nor2_1
X_26220_ _02163_ _04359_ VPWR VGND _06486_ sg13g2_nor2_1
X_26221_ _04356_ _06485_ _06486_ _04362_ VPWR VGND 
+ _06487_
+ sg13g2_a22oi_1
X_26222_ _02140_ _03822_ VPWR VGND _06488_ sg13g2_nand2b_1
X_26223_ _04651_ _02163_ _06488_ VPWR VGND _06489_ sg13g2_o21ai_1
X_26224_ _04364_ _06489_ _03740_ VPWR VGND _06490_ sg13g2_a21oi_1
X_26225_ _04355_ _06487_ _06490_ VPWR VGND _06491_ sg13g2_a21oi_1
X_26226_ _00127_ _04353_ _04354_ _02194_ _06491_ VPWR 
+ VGND
+ _06492_ sg13g2_a221oi_1
X_26227_ _00125_ _03732_ VPWR VGND _06493_ sg13g2_nand2_1
X_26228_ \atbs_core_0.spike_memory_0.n2409_o[5]\ _04373_ _06493_ VPWR VGND _06494_ sg13g2_o21ai_1
X_26229_ _04379_ _02623_ VPWR VGND _06495_ sg13g2_nor2_1
X_26230_ _02645_ _04381_ VPWR VGND _06496_ sg13g2_nor2_1
X_26231_ _04511_ _06495_ _06496_ _04384_ VPWR VGND 
+ _06497_
+ sg13g2_a22oi_1
X_26232_ _02623_ _04268_ VPWR VGND _06498_ sg13g2_nand2b_1
X_26233_ _04383_ _02645_ _06498_ VPWR VGND _06499_ sg13g2_o21ai_1
X_26234_ _04517_ _06499_ _04521_ VPWR VGND _06500_ sg13g2_a21oi_1
X_26235_ _04377_ _06497_ _06500_ VPWR VGND _06501_ sg13g2_a21oi_1
X_26236_ _12078_ _06494_ _06501_ VPWR VGND _06502_ sg13g2_nor3_1
X_26237_ _03717_ _06484_ _06492_ _04371_ _06502_ VPWR 
+ VGND
+ _06503_ sg13g2_a221oi_1
X_26238_ \atbs_core_0.spike_memory_0.n2436_q[1202]\ _03776_ VPWR VGND _06504_ sg13g2_nor2_1
X_26239_ \atbs_core_0.spike_memory_0.n2418_o[5]\ _03806_ VPWR VGND _06505_ sg13g2_nor2_1
X_26240_ _03855_ _12635_ VPWR VGND _06506_ sg13g2_nor2_1
X_26241_ _12660_ _03951_ VPWR VGND _06507_ sg13g2_nor2_1
X_26242_ _04047_ _06506_ _06507_ _04052_ VPWR VGND 
+ _06508_
+ sg13g2_a22oi_1
X_26243_ _12635_ _04054_ VPWR VGND _06509_ sg13g2_nand2b_1
X_26244_ _04051_ _12660_ _06509_ VPWR VGND _06510_ sg13g2_o21ai_1
X_26245_ _03955_ _06510_ _03868_ VPWR VGND _06511_ sg13g2_a21oi_1
X_26246_ _03993_ _06508_ _06511_ VPWR VGND _06512_ sg13g2_a21oi_1
X_26247_ _12094_ _06504_ _06505_ _06512_ VPWR VGND 
+ _06513_
+ sg13g2_nor4_1
X_26248_ \atbs_core_0.spike_memory_0.n2417_o[5]\ _04260_ VPWR VGND _06514_ sg13g2_nor2_1
X_26249_ \atbs_core_0.spike_memory_0.n2414_o[5]\ _03835_ _03780_ VPWR VGND _06515_ sg13g2_o21ai_1
X_26250_ _04089_ _12578_ VPWR VGND _06516_ sg13g2_nor2_1
X_26251_ _12601_ _04086_ VPWR VGND _06517_ sg13g2_nor2_1
X_26252_ _04082_ _06516_ _06517_ _04090_ VPWR VGND 
+ _06518_
+ sg13g2_a22oi_1
X_26253_ _12578_ _04094_ VPWR VGND _06519_ sg13g2_nand2b_1
X_26254_ _04413_ _12601_ _06519_ VPWR VGND _06520_ sg13g2_o21ai_1
X_26255_ _04092_ _06520_ _04839_ VPWR VGND _06521_ sg13g2_a21oi_1
X_26256_ _04081_ _06518_ _06521_ VPWR VGND _06522_ sg13g2_a21oi_1
X_26257_ _06514_ _06515_ _06522_ VPWR VGND _06523_ sg13g2_nor3_1
X_26258_ \atbs_core_0.spike_memory_0.n2413_o[5]\ _03803_ VPWR VGND _06524_ sg13g2_nor2_1
X_26259_ \atbs_core_0.spike_memory_0.n2410_o[5]\ _04102_ VPWR VGND _06525_ sg13g2_nor2_1
X_26260_ _03989_ _12522_ VPWR VGND _06526_ sg13g2_nor2_1
X_26261_ _12546_ _03851_ VPWR VGND _06527_ sg13g2_nor2_1
X_26262_ _04280_ _06526_ _06527_ _04283_ VPWR VGND 
+ _06528_
+ sg13g2_a22oi_1
X_26263_ _12522_ _03982_ VPWR VGND _06529_ sg13g2_nand2b_1
X_26264_ _03847_ _12546_ _06529_ VPWR VGND _06530_ sg13g2_o21ai_1
X_26265_ _03860_ _06530_ _04287_ VPWR VGND _06531_ sg13g2_a21oi_1
X_26266_ _04392_ _06528_ _06531_ VPWR VGND _06532_ sg13g2_a21oi_1
X_26267_ _03800_ _06524_ _06525_ _06532_ VPWR VGND 
+ _06533_
+ sg13g2_nor4_1
X_26268_ _06513_ _06523_ _06533_ VPWR VGND _06534_ sg13g2_nor3_1
X_26269_ \atbs_core_0.spike_memory_0.n2385_o[5]\ _03970_ VPWR VGND _06535_ sg13g2_nand2b_1
X_26270_ \atbs_core_0.spike_memory_0.n2382_o[5]\ _04292_ _06535_ VPWR VGND _06536_ sg13g2_o21ai_1
X_26271_ _04011_ _02293_ VPWR VGND _06537_ sg13g2_nor2_1
X_26272_ _02315_ _04085_ VPWR VGND _06538_ sg13g2_nor2_1
X_26273_ _03750_ _06537_ _06538_ _03989_ VPWR VGND 
+ _06539_
+ sg13g2_a22oi_1
X_26274_ _02293_ _04093_ VPWR VGND _06540_ sg13g2_nand2b_1
X_26275_ _04088_ _02315_ _06540_ VPWR VGND _06541_ sg13g2_o21ai_1
X_26276_ _03859_ _06541_ _04097_ VPWR VGND _06542_ sg13g2_a21oi_1
X_26277_ _03768_ _06539_ _06542_ VPWR VGND _06543_ sg13g2_a21oi_1
X_26278_ _06536_ _06543_ VPWR VGND _06544_ sg13g2_or2_1
X_26279_ \atbs_core_0.spike_memory_0.n2381_o[5]\ _12084_ VPWR VGND _06545_ sg13g2_nor2_1
X_26280_ \atbs_core_0.spike_memory_0.n2378_o[5]\ _03999_ VPWR VGND _06546_ sg13g2_nor2_1
X_26281_ _03890_ _02237_ VPWR VGND _06547_ sg13g2_nor2_1
X_26282_ _02260_ _03741_ VPWR VGND _06548_ sg13g2_nor2_1
X_26283_ _03850_ _06547_ _06548_ _03791_ VPWR VGND 
+ _06549_
+ sg13g2_a22oi_1
X_26284_ _02237_ _02709_ VPWR VGND _06550_ sg13g2_nand2b_1
X_26285_ _03890_ _02260_ _06550_ VPWR VGND _06551_ sg13g2_o21ai_1
X_26286_ _03730_ _06551_ _02698_ VPWR VGND _06552_ sg13g2_a21oi_1
X_26287_ _03867_ _06549_ _06552_ VPWR VGND _06553_ sg13g2_a21oi_1
X_26288_ _03726_ _06545_ _06546_ _06553_ VPWR VGND 
+ _06554_
+ sg13g2_nor4_1
X_26289_ \atbs_core_0.spike_memory_0.n2389_o[5]\ _04442_ VPWR VGND _06555_ sg13g2_nor2_1
X_26290_ \atbs_core_0.spike_memory_0.n2386_o[5]\ _03999_ VPWR VGND _06556_ sg13g2_nor2_1
X_26291_ _04455_ _02347_ VPWR VGND _06557_ sg13g2_nor2_1
X_26292_ _02371_ _03741_ VPWR VGND _06558_ sg13g2_nor2_1
X_26293_ _04085_ _06557_ _06558_ _03791_ VPWR VGND 
+ _06559_
+ sg13g2_a22oi_1
X_26294_ _02347_ _03845_ VPWR VGND _06560_ sg13g2_nand2b_1
X_26295_ _03890_ _02371_ _06560_ VPWR VGND _06561_ sg13g2_o21ai_1
X_26296_ _03730_ _06561_ _03809_ VPWR VGND _06562_ sg13g2_a21oi_1
X_26297_ _04068_ _06559_ _06562_ VPWR VGND _06563_ sg13g2_a21oi_1
X_26298_ _07555_ _06555_ _06556_ _06563_ VPWR VGND 
+ _06564_
+ sg13g2_nor4_1
X_26299_ _06554_ _06564_ _12090_ VPWR VGND _06565_ sg13g2_o21ai_1
X_26300_ _04276_ _06544_ _06565_ VPWR VGND _06566_ sg13g2_o21ai_1
X_26301_ \atbs_core_0.spike_memory_0.n2401_o[5]\ _03970_ VPWR VGND _06567_ sg13g2_nand2b_1
X_26302_ \atbs_core_0.spike_memory_0.n2398_o[5]\ _04078_ _06567_ VPWR VGND _06568_ sg13g2_o21ai_1
X_26303_ _03891_ _02529_ VPWR VGND _06569_ sg13g2_nor2_1
X_26304_ _02550_ _04107_ VPWR VGND _06570_ sg13g2_nor2_1
X_26305_ _03818_ _06569_ _06570_ _04346_ VPWR VGND 
+ _06571_
+ sg13g2_a22oi_1
X_26306_ _02529_ _02710_ VPWR VGND _06572_ sg13g2_nand2b_1
X_26307_ _03763_ _02550_ _06572_ VPWR VGND _06573_ sg13g2_o21ai_1
X_26308_ _03986_ _06573_ _02699_ VPWR VGND _06574_ sg13g2_a21oi_1
X_26309_ _03830_ _06571_ _06574_ VPWR VGND _06575_ sg13g2_a21oi_1
X_26310_ _06568_ _06575_ VPWR VGND _06576_ sg13g2_or2_1
X_26311_ \atbs_core_0.spike_memory_0.n2397_o[5]\ _04442_ VPWR VGND _06577_ sg13g2_nor2_1
X_26312_ \atbs_core_0.spike_memory_0.n2394_o[5]\ _03999_ VPWR VGND _06578_ sg13g2_nor2_1
X_26313_ _03862_ _02480_ VPWR VGND _06579_ sg13g2_nor2_1
X_26314_ _02502_ _03749_ VPWR VGND _06580_ sg13g2_nor2_1
X_26315_ _04085_ _06579_ _06580_ _04480_ VPWR VGND 
+ _06581_
+ sg13g2_a22oi_1
X_26316_ _02480_ _03845_ VPWR VGND _06582_ sg13g2_nand2b_1
X_26317_ _03862_ _02502_ _06582_ VPWR VGND _06583_ sg13g2_o21ai_1
X_26318_ _04009_ _06583_ _03809_ VPWR VGND _06584_ sg13g2_a21oi_1
X_26319_ _04097_ _06581_ _06584_ VPWR VGND _06585_ sg13g2_a21oi_1
X_26320_ _03726_ _06577_ _06578_ _06585_ VPWR VGND 
+ _06586_
+ sg13g2_nor4_1
X_26321_ \atbs_core_0.spike_memory_0.n2405_o[5]\ _04442_ VPWR VGND _06587_ sg13g2_nor2_1
X_26322_ \atbs_core_0.spike_memory_0.n2402_o[5]\ _03778_ VPWR VGND _06588_ sg13g2_nor2_1
X_26323_ _04093_ _02576_ VPWR VGND _06589_ sg13g2_nor2_1
X_26324_ _02597_ _03749_ VPWR VGND _06590_ sg13g2_nor2_1
X_26325_ _04107_ _06589_ _06590_ _03982_ VPWR VGND 
+ _06591_
+ sg13g2_a22oi_1
X_26326_ _02576_ _03762_ VPWR VGND _06592_ sg13g2_nand2b_1
X_26327_ _03981_ _02597_ _06592_ VPWR VGND _06593_ sg13g2_o21ai_1
X_26328_ _04009_ _06593_ _03809_ VPWR VGND _06594_ sg13g2_a21oi_1
X_26329_ _04097_ _06591_ _06594_ VPWR VGND _06595_ sg13g2_a21oi_1
X_26330_ _07555_ _06587_ _06588_ _06595_ VPWR VGND 
+ _06596_
+ sg13g2_nor4_1
X_26331_ _06586_ _06596_ _12090_ VPWR VGND _06597_ sg13g2_o21ai_1
X_26332_ _04276_ _06576_ _06597_ VPWR VGND _06598_ sg13g2_o21ai_1
X_26333_ _07547_ _06566_ _06598_ _03717_ VPWR VGND 
+ _06599_
+ sg13g2_a22oi_1
X_26334_ _12079_ _06534_ _06599_ VPWR VGND _06600_ sg13g2_o21ai_1
X_26335_ _04336_ _06600_ VPWR VGND _06601_ sg13g2_nor2_1
X_26336_ _04336_ _06503_ _06601_ VPWR VGND _06602_ sg13g2_a21oi_1
X_26337_ \atbs_core_0.spike_memory_0.n2361_o[5]\ _04373_ VPWR VGND _06603_ sg13g2_nor2_1
X_26338_ \atbs_core_0.spike_memory_0.n2358_o[5]\ _04606_ VPWR VGND _06604_ sg13g2_nor2_1
X_26339_ _04513_ _02082_ VPWR VGND _06605_ sg13g2_nor2_1
X_26340_ _02277_ _04716_ VPWR VGND _06606_ sg13g2_nor2_1
X_26341_ _04511_ _06605_ _06606_ _04613_ VPWR VGND 
+ _06607_
+ sg13g2_a22oi_1
X_26342_ _02082_ _04518_ VPWR VGND _06608_ sg13g2_nand2b_1
X_26343_ _03984_ _02277_ _06608_ VPWR VGND _06609_ sg13g2_o21ai_1
X_26344_ _04517_ _06609_ _04521_ VPWR VGND _06610_ sg13g2_a21oi_1
X_26345_ _04608_ _06607_ _06610_ VPWR VGND _06611_ sg13g2_a21oi_1
X_26346_ _04505_ _06603_ _06604_ _06611_ VPWR VGND 
+ _06612_
+ sg13g2_nor4_1
X_26347_ \atbs_core_0.spike_memory_0.n2369_o[5]\ _04525_ VPWR VGND _06613_ sg13g2_nor2_1
X_26348_ \atbs_core_0.spike_memory_0.n2366_o[5]\ _04549_ VPWR VGND _06614_ sg13g2_nor2_1
X_26349_ _04553_ _02031_ VPWR VGND _06615_ sg13g2_nor2_1
X_26350_ _02052_ _04533_ VPWR VGND _06616_ sg13g2_nor2_1
X_26351_ _04531_ _06615_ _06616_ _04557_ VPWR VGND 
+ _06617_
+ sg13g2_a22oi_1
X_26352_ _02031_ _04559_ VPWR VGND _06618_ sg13g2_nand2b_1
X_26353_ _04539_ _02052_ _06618_ VPWR VGND _06619_ sg13g2_o21ai_1
X_26354_ _04538_ _06619_ _04562_ VPWR VGND _06620_ sg13g2_a21oi_1
X_26355_ _04551_ _06617_ _06620_ VPWR VGND _06621_ sg13g2_a21oi_1
X_26356_ _04604_ _06613_ _06614_ _06621_ VPWR VGND 
+ _06622_
+ sg13g2_nor4_1
X_26357_ _03925_ _06612_ _06622_ VPWR VGND _06623_ sg13g2_nor3_1
X_26358_ \atbs_core_0.spike_memory_0.n2365_o[5]\ _04506_ VPWR VGND _06624_ sg13g2_nor2_1
X_26359_ \atbs_core_0.spike_memory_0.n2362_o[5]\ _04508_ VPWR VGND _06625_ sg13g2_nor2_1
X_26360_ _04535_ _12519_ VPWR VGND _06626_ sg13g2_nor2_1
X_26361_ _12678_ _04555_ VPWR VGND _06627_ sg13g2_nor2_1
X_26362_ _04378_ _06626_ _06627_ _04384_ VPWR VGND 
+ _06628_
+ sg13g2_a22oi_1
X_26363_ _12519_ _05544_ VPWR VGND _06629_ sg13g2_nand2b_1
X_26364_ _03755_ _12678_ _06629_ VPWR VGND _06630_ sg13g2_o21ai_1
X_26365_ _04388_ _06630_ _04393_ VPWR VGND _06631_ sg13g2_a21oi_1
X_26366_ _04377_ _06628_ _06631_ VPWR VGND _06632_ sg13g2_a21oi_1
X_26367_ _03968_ _06624_ _06625_ _06632_ VPWR VGND 
+ _06633_
+ sg13g2_nor4_1
X_26368_ \atbs_core_0.spike_memory_0.n2373_o[5]\ _12088_ VPWR VGND _06634_ sg13g2_nor2_1
X_26369_ \atbs_core_0.spike_memory_0.n2370_o[5]\ _04528_ VPWR VGND _06635_ sg13g2_nor2_1
X_26370_ _03934_ _02085_ VPWR VGND _06636_ sg13g2_nor2_1
X_26371_ _02108_ _04570_ VPWR VGND _06637_ sg13g2_nor2_1
X_26372_ _04568_ _06636_ _06637_ _04536_ VPWR VGND 
+ _06638_
+ sg13g2_a22oi_1
X_26373_ _02085_ _04361_ VPWR VGND _06639_ sg13g2_nand2b_1
X_26374_ _04574_ _02108_ _06639_ VPWR VGND _06640_ sg13g2_o21ai_1
X_26375_ _04573_ _06640_ _04542_ VPWR VGND _06641_ sg13g2_a21oi_1
X_26376_ _04530_ _06638_ _06641_ VPWR VGND _06642_ sg13g2_a21oi_1
X_26377_ _04126_ _06634_ _06635_ _06642_ VPWR VGND 
+ _06643_
+ sg13g2_nor4_1
X_26378_ _04547_ _06633_ _06643_ VPWR VGND _06644_ sg13g2_nor3_1
X_26379_ _07549_ _06623_ _06644_ VPWR VGND _06645_ sg13g2_nor3_1
X_26380_ _04503_ _06602_ _06645_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[5]\ sg13g2_a21o_1
X_26381_ _03761_ _02141_ VPWR VGND _06646_ sg13g2_nor2_1
X_26382_ _02164_ _03751_ VPWR VGND _06647_ sg13g2_nor2_1
X_26383_ _04510_ _06646_ _06647_ _04513_ VPWR VGND 
+ _06648_
+ sg13g2_a22oi_1
X_26384_ _02141_ _04111_ VPWR VGND _06649_ sg13g2_nand2b_1
X_26385_ _03978_ _02164_ _06649_ VPWR VGND _06650_ sg13g2_o21ai_1
X_26386_ _04387_ _06650_ _03840_ VPWR VGND _06651_ sg13g2_a21oi_1
X_26387_ _04376_ _06648_ _06651_ VPWR VGND _06652_ sg13g2_a21oi_1
X_26388_ _00130_ _03969_ _03972_ _02196_ _06652_ VPWR 
+ VGND
+ _06653_ sg13g2_a221oi_1
X_26389_ \atbs_core_0.spike_memory_0.n2385_o[6]\ _12086_ VPWR VGND _06654_ sg13g2_nor2_1
X_26390_ \atbs_core_0.spike_memory_0.n2382_o[6]\ _04771_ _03780_ VPWR VGND _06655_ sg13g2_o21ai_1
X_26391_ _03787_ _02294_ VPWR VGND _06656_ sg13g2_nor2_1
X_26392_ _02317_ _03750_ VPWR VGND _06657_ sg13g2_nor2_1
X_26393_ _03743_ _06656_ _06657_ _03754_ VPWR VGND 
+ _06658_
+ sg13g2_a22oi_1
X_26394_ _02294_ _03763_ VPWR VGND _06659_ sg13g2_nand2b_1
X_26395_ _03753_ _02317_ _06659_ VPWR VGND _06660_ sg13g2_o21ai_1
X_26396_ _03758_ _06660_ _04294_ VPWR VGND _06661_ sg13g2_a21oi_1
X_26397_ _03739_ _06658_ _06661_ VPWR VGND _06662_ sg13g2_a21oi_1
X_26398_ _06654_ _06655_ _06662_ VPWR VGND _06663_ sg13g2_or3_1
X_26399_ _03775_ _06663_ VPWR VGND _06664_ sg13g2_nand2_1
X_26400_ _03729_ _06653_ _06664_ VPWR VGND _06665_ sg13g2_o21ai_1
X_26401_ \atbs_core_0.spike_memory_0.n2381_o[6]\ _03944_ VPWR VGND _06666_ sg13g2_nor2_1
X_26402_ \atbs_core_0.spike_memory_0.n2378_o[6]\ _03807_ VPWR VGND _06667_ sg13g2_nor2_1
X_26403_ _03826_ _02238_ VPWR VGND _06668_ sg13g2_nor2_1
X_26404_ _02262_ _04152_ VPWR VGND _06669_ sg13g2_nor2_1
X_26405_ _04150_ _06668_ _06669_ _04154_ VPWR VGND 
+ _06670_
+ sg13g2_a22oi_1
X_26406_ _02238_ _05745_ VPWR VGND _06671_ sg13g2_nand2b_1
X_26407_ _05753_ _02262_ _06671_ VPWR VGND _06672_ sg13g2_o21ai_1
X_26408_ _03936_ _06672_ _04158_ VPWR VGND _06673_ sg13g2_a21oi_1
X_26409_ _04149_ _06670_ _06673_ VPWR VGND _06674_ sg13g2_a21oi_1
X_26410_ _06666_ _06667_ _06674_ VPWR VGND _06675_ sg13g2_nor3_1
X_26411_ \atbs_core_0.spike_memory_0.n2389_o[6]\ _03971_ VPWR VGND _06676_ sg13g2_nand2b_1
X_26412_ \atbs_core_0.spike_memory_0.n2386_o[6]\ _03836_ _06676_ VPWR VGND _06677_ sg13g2_o21ai_1
X_26413_ _03856_ _02348_ VPWR VGND _06678_ sg13g2_nor2_1
X_26414_ _02372_ _03952_ VPWR VGND _06679_ sg13g2_nor2_1
X_26415_ _03844_ _06678_ _06679_ _03857_ VPWR VGND 
+ _06680_
+ sg13g2_a22oi_1
X_26416_ _02348_ _04167_ VPWR VGND _06681_ sg13g2_nand2b_1
X_26417_ _03949_ _02372_ _06681_ VPWR VGND _06682_ sg13g2_o21ai_1
X_26418_ _03956_ _06682_ _04317_ VPWR VGND _06683_ sg13g2_a21oi_1
X_26419_ _03948_ _06680_ _06683_ VPWR VGND _06684_ sg13g2_a21oi_1
X_26420_ _06677_ _06684_ _03775_ VPWR VGND _06685_ sg13g2_o21ai_1
X_26421_ _03801_ _06675_ _06685_ VPWR VGND _06686_ sg13g2_o21ai_1
X_26422_ _03725_ _06665_ _06686_ _06663_ VPWR VGND 
+ _06687_
+ sg13g2_a22oi_1
X_26423_ _05850_ _02625_ VPWR VGND _06688_ sg13g2_nor2_1
X_26424_ _02646_ _03813_ VPWR VGND _06689_ sg13g2_nor2_1
X_26425_ _04587_ _06688_ _06689_ _04610_ VPWR VGND 
+ _06690_
+ sg13g2_a22oi_1
X_26426_ _02625_ _05533_ VPWR VGND _06691_ sg13g2_nand2b_1
X_26427_ _04589_ _02646_ _06691_ VPWR VGND _06692_ sg13g2_o21ai_1
X_26428_ _03987_ _06692_ _03811_ VPWR VGND _06693_ sg13g2_a21oi_1
X_26429_ _03974_ _06690_ _06693_ VPWR VGND _06694_ sg13g2_a21oi_1
X_26430_ _00128_ _03969_ _03972_ _02671_ _06694_ VPWR 
+ VGND
+ _06695_ sg13g2_a221oi_1
X_26431_ \atbs_core_0.spike_memory_0.n2417_o[6]\ _03876_ VPWR VGND _06696_ sg13g2_nor2_1
X_26432_ \atbs_core_0.spike_memory_0.n2414_o[6]\ _04229_ _03722_ VPWR VGND _06697_ sg13g2_o21ai_1
X_26433_ _03977_ _12579_ VPWR VGND _06698_ sg13g2_nor2_1
X_26434_ _12602_ _03842_ VPWR VGND _06699_ sg13g2_nor2_1
X_26435_ _03975_ _06698_ _06699_ _05850_ VPWR VGND 
+ _06700_
+ sg13g2_a22oi_1
X_26436_ _12579_ _04088_ VPWR VGND _06701_ sg13g2_nand2b_1
X_26437_ _04094_ _12602_ _06701_ VPWR VGND _06702_ sg13g2_o21ai_1
X_26438_ _04010_ _06702_ _03992_ VPWR VGND _06703_ sg13g2_a21oi_1
X_26439_ _04002_ _06700_ _06703_ VPWR VGND _06704_ sg13g2_a21oi_1
X_26440_ _06696_ _06697_ _06704_ VPWR VGND _06705_ sg13g2_or3_1
X_26441_ _03926_ _06705_ VPWR VGND _06706_ sg13g2_nand2_1
X_26442_ _03968_ _06695_ _06706_ VPWR VGND _06707_ sg13g2_o21ai_1
X_26443_ \atbs_core_0.spike_memory_0.n2413_o[6]\ _03877_ VPWR VGND _06708_ sg13g2_nor2_1
X_26444_ \atbs_core_0.spike_memory_0.n2410_o[6]\ _04527_ VPWR VGND _06709_ sg13g2_nor2_1
X_26445_ _03886_ _12523_ VPWR VGND _06710_ sg13g2_nor2_1
X_26446_ _12547_ _04082_ VPWR VGND _06711_ sg13g2_nor2_1
X_26447_ _03744_ _06710_ _06711_ _04539_ VPWR VGND 
+ _06712_
+ sg13g2_a22oi_1
X_26448_ _12523_ _04105_ VPWR VGND _06713_ sg13g2_nand2b_1
X_26449_ _03747_ _12547_ _06713_ VPWR VGND _06714_ sg13g2_o21ai_1
X_26450_ _03759_ _06714_ _03769_ VPWR VGND _06715_ sg13g2_a21oi_1
X_26451_ _03740_ _06712_ _06715_ VPWR VGND _06716_ sg13g2_a21oi_1
X_26452_ _06708_ _06709_ _06716_ VPWR VGND _06717_ sg13g2_nor3_1
X_26453_ \atbs_core_0.spike_memory_0.n2436_q[1203]\ _03971_ VPWR VGND _06718_ sg13g2_nand2b_1
X_26454_ \atbs_core_0.spike_memory_0.n2418_o[6]\ _04032_ _06718_ VPWR VGND _06719_ sg13g2_o21ai_1
X_26455_ _03826_ _12636_ VPWR VGND _06720_ sg13g2_nor2_1
X_26456_ _12661_ _03932_ VPWR VGND _06721_ sg13g2_nor2_1
X_26457_ _03929_ _06720_ _06721_ _03934_ VPWR VGND 
+ _06722_
+ sg13g2_a22oi_1
X_26458_ _12636_ _03937_ VPWR VGND _06723_ sg13g2_nand2b_1
X_26459_ _02712_ _12661_ _06723_ VPWR VGND _06724_ sg13g2_o21ai_1
X_26460_ _03936_ _06724_ _04158_ VPWR VGND _06725_ sg13g2_a21oi_1
X_26461_ _02701_ _06722_ _06725_ VPWR VGND _06726_ sg13g2_a21oi_1
X_26462_ _06719_ _06726_ _03997_ VPWR VGND _06727_ sg13g2_o21ai_1
X_26463_ _04074_ _06717_ _06727_ VPWR VGND _06728_ sg13g2_o21ai_1
X_26464_ _03967_ _06707_ _06728_ _06705_ _04045_ VPWR 
+ VGND
+ _06729_ sg13g2_a221oi_1
X_26465_ _03721_ _06687_ _06729_ VPWR VGND _06730_ sg13g2_a21oi_1
X_26466_ \atbs_core_0.spike_memory_0.n2369_o[6]\ _03803_ VPWR VGND _06731_ sg13g2_nor2_1
X_26467_ \atbs_core_0.spike_memory_0.n2366_o[6]\ _03806_ VPWR VGND _06732_ sg13g2_nor2_1
X_26468_ _03815_ _02032_ VPWR VGND _06733_ sg13g2_nor2_1
X_26469_ _02053_ _03951_ VPWR VGND _06734_ sg13g2_nor2_1
X_26470_ _03813_ _06733_ _06734_ _03907_ VPWR VGND 
+ _06735_
+ sg13g2_a22oi_1
X_26471_ _02032_ _03915_ VPWR VGND _06736_ sg13g2_nand2b_1
X_26472_ _03821_ _02053_ _06736_ VPWR VGND _06737_ sg13g2_o21ai_1
X_26473_ _03790_ _06737_ _03830_ VPWR VGND _06738_ sg13g2_a21oi_1
X_26474_ _03811_ _06735_ _06738_ VPWR VGND _06739_ sg13g2_a21oi_1
X_26475_ _06731_ _06732_ _06739_ VPWR VGND _06740_ sg13g2_nor3_1
X_26476_ \atbs_core_0.spike_memory_0.n2361_o[6]\ _03776_ VPWR VGND _06741_ sg13g2_nor2_1
X_26477_ \atbs_core_0.spike_memory_0.n2358_o[6]\ _05540_ VPWR VGND _06742_ sg13g2_nor2_1
X_26478_ _03855_ _02094_ VPWR VGND _06743_ sg13g2_nor2_1
X_26479_ _02280_ _03951_ VPWR VGND _06744_ sg13g2_nor2_1
X_26480_ _03843_ _06743_ _06744_ _03949_ VPWR VGND 
+ _06745_
+ sg13g2_a22oi_1
X_26481_ _02094_ _04054_ VPWR VGND _06746_ sg13g2_nand2b_1
X_26482_ _04051_ _02280_ _06746_ VPWR VGND _06747_ sg13g2_o21ai_1
X_26483_ _03955_ _06747_ _03868_ VPWR VGND _06748_ sg13g2_a21oi_1
X_26484_ _03993_ _06745_ _06748_ VPWR VGND _06749_ sg13g2_a21oi_1
X_26485_ _04244_ _06741_ _06742_ _06749_ VPWR VGND 
+ _06750_
+ sg13g2_nor4_1
X_26486_ _03926_ _06740_ _06750_ VPWR VGND _06751_ sg13g2_a21oi_1
X_26487_ \atbs_core_0.spike_memory_0.n2365_o[6]\ _03776_ VPWR VGND _06752_ sg13g2_nor2_1
X_26488_ \atbs_core_0.spike_memory_0.n2362_o[6]\ _03806_ VPWR VGND _06753_ sg13g2_nor2_1
X_26489_ _04051_ _12532_ VPWR VGND _06754_ sg13g2_nor2_1
X_26490_ _12681_ _03951_ VPWR VGND _06755_ sg13g2_nor2_1
X_26491_ _04047_ _06754_ _06755_ _03957_ VPWR VGND 
+ _06756_
+ sg13g2_a22oi_1
X_26492_ _12532_ _04054_ VPWR VGND _06757_ sg13g2_nand2b_1
X_26493_ _03815_ _12681_ _06757_ VPWR VGND _06758_ sg13g2_o21ai_1
X_26494_ _03955_ _06758_ _03830_ VPWR VGND _06759_ sg13g2_a21oi_1
X_26495_ _03993_ _06756_ _06759_ VPWR VGND _06760_ sg13g2_a21oi_1
X_26496_ _03727_ _06752_ _06753_ _06760_ VPWR VGND 
+ _06761_
+ sg13g2_nor4_1
X_26497_ \atbs_core_0.spike_memory_0.n2373_o[6]\ _03803_ VPWR VGND _06762_ sg13g2_nor2_1
X_26498_ \atbs_core_0.spike_memory_0.n2370_o[6]\ _04102_ VPWR VGND _06763_ sg13g2_nor2_1
X_26499_ _03847_ _02086_ VPWR VGND _06764_ sg13g2_nor2_1
X_26500_ _02110_ _03851_ VPWR VGND _06765_ sg13g2_nor2_1
X_26501_ _03843_ _06764_ _06765_ _04708_ VPWR VGND 
+ _06766_
+ sg13g2_a22oi_1
X_26502_ _02086_ _03982_ VPWR VGND _06767_ sg13g2_nand2b_1
X_26503_ _04597_ _02110_ _06767_ VPWR VGND _06768_ sg13g2_o21ai_1
X_26504_ _03860_ _06768_ _04287_ VPWR VGND _06769_ sg13g2_a21oi_1
X_26505_ _03840_ _06766_ _06769_ VPWR VGND _06770_ sg13g2_a21oi_1
X_26506_ _03899_ _06762_ _06763_ _06770_ VPWR VGND 
+ _06771_
+ sg13g2_nor4_1
X_26507_ _03966_ _06761_ _06771_ VPWR VGND _06772_ sg13g2_nor3_1
X_26508_ _03724_ _06751_ _06772_ VPWR VGND _06773_ sg13g2_a21oi_1
X_26509_ _04045_ _06773_ VPWR VGND _06774_ sg13g2_and2_1
X_26510_ _05850_ _02397_ VPWR VGND _06775_ sg13g2_nor2_1
X_26511_ _02416_ _04047_ VPWR VGND _06776_ sg13g2_nor2_1
X_26512_ _04587_ _06775_ _06776_ _03984_ VPWR VGND 
+ _06777_
+ sg13g2_a22oi_1
X_26513_ _02397_ _03989_ VPWR VGND _06778_ sg13g2_nand2b_1
X_26514_ _03983_ _02416_ _06778_ VPWR VGND _06779_ sg13g2_o21ai_1
X_26515_ _03987_ _06779_ _03811_ VPWR VGND _06780_ sg13g2_a21oi_1
X_26516_ _03974_ _06777_ _06780_ VPWR VGND _06781_ sg13g2_a21oi_1
X_26517_ _00129_ _03969_ _03972_ _02444_ _06781_ VPWR 
+ VGND
+ _06782_ sg13g2_a221oi_1
X_26518_ \atbs_core_0.spike_memory_0.n2401_o[6]\ _03876_ VPWR VGND _06783_ sg13g2_nor2_1
X_26519_ \atbs_core_0.spike_memory_0.n2398_o[6]\ _04229_ _03722_ VPWR VGND _06784_ sg13g2_o21ai_1
X_26520_ _03977_ _02530_ VPWR VGND _06785_ sg13g2_nor2_1
X_26521_ _02551_ _04062_ VPWR VGND _06786_ sg13g2_nor2_1
X_26522_ _03975_ _06785_ _06786_ _05850_ VPWR VGND 
+ _06787_
+ sg13g2_a22oi_1
X_26523_ _02530_ _04011_ VPWR VGND _06788_ sg13g2_nand2b_1
X_26524_ _04254_ _02551_ _06788_ VPWR VGND _06789_ sg13g2_o21ai_1
X_26525_ _04010_ _06789_ _03992_ VPWR VGND _06790_ sg13g2_a21oi_1
X_26526_ _04002_ _06787_ _06790_ VPWR VGND _06791_ sg13g2_a21oi_1
X_26527_ _06783_ _06784_ _06791_ VPWR VGND _06792_ sg13g2_or3_1
X_26528_ _03997_ _06792_ VPWR VGND _06793_ sg13g2_nand2_1
X_26529_ _03968_ _06782_ _06793_ VPWR VGND _06794_ sg13g2_o21ai_1
X_26530_ \atbs_core_0.spike_memory_0.n2397_o[6]\ _12087_ VPWR VGND _06795_ sg13g2_nor2_1
X_26531_ \atbs_core_0.spike_memory_0.n2394_o[6]\ _04527_ VPWR VGND _06796_ sg13g2_nor2_1
X_26532_ _03886_ _02481_ VPWR VGND _06797_ sg13g2_nor2_1
X_26533_ _02503_ _04023_ VPWR VGND _06798_ sg13g2_nor2_1
X_26534_ _04359_ _06797_ _06798_ _04535_ VPWR VGND 
+ _06799_
+ sg13g2_a22oi_1
X_26535_ _02481_ _04105_ VPWR VGND _06800_ sg13g2_nand2b_1
X_26536_ _03788_ _02503_ _06800_ VPWR VGND _06801_ sg13g2_o21ai_1
X_26537_ _03759_ _06801_ _03769_ VPWR VGND _06802_ sg13g2_a21oi_1
X_26538_ _04021_ _06799_ _06802_ VPWR VGND _06803_ sg13g2_a21oi_1
X_26539_ _06795_ _06796_ _06803_ VPWR VGND _06804_ sg13g2_nor3_1
X_26540_ \atbs_core_0.spike_memory_0.n2405_o[6]\ _03971_ VPWR VGND _06805_ sg13g2_nand2b_1
X_26541_ \atbs_core_0.spike_memory_0.n2402_o[6]\ _04032_ _06805_ VPWR VGND _06806_ sg13g2_o21ai_1
X_26542_ _03826_ _02577_ VPWR VGND _06807_ sg13g2_nor2_1
X_26543_ _02598_ _04152_ VPWR VGND _06808_ sg13g2_nor2_1
X_26544_ _04150_ _06807_ _06808_ _04154_ VPWR VGND 
+ _06809_
+ sg13g2_a22oi_1
X_26545_ _02577_ _03937_ VPWR VGND _06810_ sg13g2_nand2b_1
X_26546_ _05753_ _02598_ _06810_ VPWR VGND _06811_ sg13g2_o21ai_1
X_26547_ _03936_ _06811_ _04158_ VPWR VGND _06812_ sg13g2_a21oi_1
X_26548_ _02701_ _06809_ _06812_ VPWR VGND _06813_ sg13g2_a21oi_1
X_26549_ _06806_ _06813_ _03997_ VPWR VGND _06814_ sg13g2_o21ai_1
X_26550_ _03801_ _06804_ _06814_ VPWR VGND _06815_ sg13g2_o21ai_1
X_26551_ _03967_ _06794_ _06815_ _06792_ _04045_ VPWR 
+ VGND
+ _06816_ sg13g2_a221oi_1
X_26552_ _06774_ _06816_ _03719_ VPWR VGND _06817_ sg13g2_o21ai_1
X_26553_ _03719_ _06730_ _06817_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[6]\ sg13g2_o21ai_1
X_26554_ \atbs_core_0.spike_memory_0.n2365_o[7]\ _04623_ VPWR VGND _06818_ sg13g2_nor2_1
X_26555_ \atbs_core_0.spike_memory_0.n2362_o[7]\ _04584_ VPWR VGND _06819_ sg13g2_nor2_1
X_26556_ _04590_ _12544_ VPWR VGND _06820_ sg13g2_nor2_1
X_26557_ _02007_ _03929_ VPWR VGND _06821_ sg13g2_nor2_1
X_26558_ _04588_ _06820_ _06821_ _04630_ VPWR VGND 
+ _06822_
+ sg13g2_a22oi_1
X_26559_ _12544_ _04598_ VPWR VGND _06823_ sg13g2_nand2b_1
X_26560_ _04632_ _02007_ _06823_ VPWR VGND _06824_ sg13g2_o21ai_1
X_26561_ _04596_ _06824_ _04635_ VPWR VGND _06825_ sg13g2_a21oi_1
X_26562_ _04626_ _06822_ _06825_ VPWR VGND _06826_ sg13g2_a21oi_1
X_26563_ _03872_ _06818_ _06819_ _06826_ VPWR VGND 
+ _06827_
+ sg13g2_nor4_1
X_26564_ \atbs_core_0.spike_memory_0.n2373_o[7]\ _04582_ VPWR VGND _06828_ sg13g2_nor2_1
X_26565_ \atbs_core_0.spike_memory_0.n2370_o[7]\ _04606_ VPWR VGND _06829_ sg13g2_nor2_1
X_26566_ _04610_ _02088_ VPWR VGND _06830_ sg13g2_nor2_1
X_26567_ _02111_ _03814_ VPWR VGND _06831_ sg13g2_nor2_1
X_26568_ _04609_ _06830_ _06831_ _04594_ VPWR VGND 
+ _06832_
+ sg13g2_a22oi_1
X_26569_ _02088_ _04708_ VPWR VGND _06833_ sg13g2_nand2b_1
X_26570_ _04616_ _02111_ _06833_ VPWR VGND _06834_ sg13g2_o21ai_1
X_26571_ _04615_ _06834_ _03812_ VPWR VGND _06835_ sg13g2_a21oi_1
X_26572_ _04586_ _06832_ _06835_ VPWR VGND _06836_ sg13g2_a21oi_1
X_26573_ _04219_ _06828_ _06829_ _06836_ VPWR VGND 
+ _06837_
+ sg13g2_nor4_1
X_26574_ _06827_ _06837_ _04504_ VPWR VGND _06838_ sg13g2_o21ai_1
X_26575_ \atbs_core_0.spike_memory_0.n2361_o[7]\ _04623_ VPWR VGND _06839_ sg13g2_nor2_1
X_26576_ \atbs_core_0.spike_memory_0.n2358_o[7]\ _03946_ VPWR VGND _06840_ sg13g2_nor2_1
X_26577_ _04593_ _02106_ VPWR VGND _06841_ sg13g2_nor2_1
X_26578_ _02282_ _04628_ VPWR VGND _06842_ sg13g2_nor2_1
X_26579_ _04662_ _06841_ _06842_ _04630_ VPWR VGND 
+ _06843_
+ sg13g2_a22oi_1
X_26580_ _02106_ _04052_ VPWR VGND _06844_ sg13g2_nand2b_1
X_26581_ _04357_ _02282_ _06844_ VPWR VGND _06845_ sg13g2_o21ai_1
X_26582_ _04666_ _06845_ _03880_ VPWR VGND _06846_ sg13g2_a21oi_1
X_26583_ _04626_ _06843_ _06846_ VPWR VGND _06847_ sg13g2_a21oi_1
X_26584_ _03872_ _06839_ _06840_ _06847_ VPWR VGND 
+ _06848_
+ sg13g2_nor4_1
X_26585_ \atbs_core_0.spike_memory_0.n2369_o[7]\ _04582_ VPWR VGND _06849_ sg13g2_nor2_1
X_26586_ \atbs_core_0.spike_memory_0.n2366_o[7]\ _04584_ VPWR VGND _06850_ sg13g2_nor2_1
X_26587_ _04616_ _02033_ VPWR VGND _06851_ sg13g2_nor2_1
X_26588_ _02054_ _03906_ VPWR VGND _06852_ sg13g2_nor2_1
X_26589_ _04588_ _06851_ _06852_ _04594_ VPWR VGND 
+ _06853_
+ sg13g2_a22oi_1
X_26590_ _02033_ _03856_ VPWR VGND _06854_ sg13g2_nand2b_1
X_26591_ _04590_ _02054_ _06854_ VPWR VGND _06855_ sg13g2_o21ai_1
X_26592_ _04596_ _06855_ _04149_ VPWR VGND _06856_ sg13g2_a21oi_1
X_26593_ _04586_ _06853_ _06856_ VPWR VGND _06857_ sg13g2_a21oi_1
X_26594_ _04219_ _06849_ _06850_ _06857_ VPWR VGND 
+ _06858_
+ sg13g2_nor4_1
X_26595_ _06848_ _06858_ _03725_ VPWR VGND _06859_ sg13g2_o21ai_1
X_26596_ _06838_ _06859_ VPWR VGND _06860_ sg13g2_and2_1
X_26597_ _04651_ _02398_ VPWR VGND _06861_ sg13g2_nor2_1
X_26598_ _02417_ _04510_ VPWR VGND _06862_ sg13g2_nor2_1
X_26599_ _04356_ _06861_ _06862_ _04680_ VPWR VGND 
+ _06863_
+ sg13g2_a22oi_1
X_26600_ _02398_ _04552_ VPWR VGND _06864_ sg13g2_nand2b_1
X_26601_ _04320_ _02417_ _06864_ VPWR VGND _06865_ sg13g2_o21ai_1
X_26602_ _04364_ _06865_ _04684_ VPWR VGND _06866_ sg13g2_a21oi_1
X_26603_ _04677_ _06863_ _06866_ VPWR VGND _06867_ sg13g2_a21oi_1
X_26604_ _00132_ _04675_ _04676_ _02446_ _06867_ VPWR 
+ VGND
+ _06868_ sg13g2_a221oi_1
X_26605_ _04632_ _02626_ VPWR VGND _06869_ sg13g2_nor2_1
X_26606_ _02647_ _03881_ VPWR VGND _06870_ sg13g2_nor2_1
X_26607_ _04662_ _06869_ _06870_ _04362_ VPWR VGND 
+ _06871_
+ sg13g2_a22oi_1
X_26608_ _02626_ _03957_ VPWR VGND _06872_ sg13g2_nand2b_1
X_26609_ _04365_ _02647_ _06872_ VPWR VGND _06873_ sg13g2_o21ai_1
X_26610_ _04666_ _06873_ _04021_ VPWR VGND _06874_ sg13g2_a21oi_1
X_26611_ _04355_ _06871_ _06874_ VPWR VGND _06875_ sg13g2_a21oi_1
X_26612_ _00131_ _04353_ _04354_ _02673_ _06875_ VPWR 
+ VGND
+ _06876_ sg13g2_a221oi_1
X_26613_ _04337_ _06868_ _06876_ _04673_ VPWR VGND 
+ _06877_
+ sg13g2_a22oi_1
X_26614_ _04361_ _02143_ VPWR VGND _06878_ sg13g2_nor2_1
X_26615_ _02165_ _03976_ VPWR VGND _06879_ sg13g2_nor2_1
X_26616_ _04339_ _06878_ _06879_ _04680_ VPWR VGND 
+ _06880_
+ sg13g2_a22oi_1
X_26617_ _02143_ _04552_ VPWR VGND _06881_ sg13g2_nand2b_1
X_26618_ _04340_ _02165_ _06881_ VPWR VGND _06882_ sg13g2_o21ai_1
X_26619_ _04345_ _06882_ _04684_ VPWR VGND _06883_ sg13g2_a21oi_1
X_26620_ _04677_ _06880_ _06883_ VPWR VGND _06884_ sg13g2_a21oi_1
X_26621_ _00133_ _04675_ _04676_ _02198_ _06884_ VPWR 
+ VGND
+ _06885_ sg13g2_a221oi_1
X_26622_ _04371_ _06885_ _04688_ VPWR VGND _06886_ sg13g2_a21oi_1
X_26623_ _06877_ _06886_ VPWR VGND _06887_ sg13g2_nand2_1
X_26624_ \atbs_core_0.spike_memory_0.n2413_o[7]\ _03901_ VPWR VGND _06888_ sg13g2_nor2_1
X_26625_ \atbs_core_0.spike_memory_0.n2410_o[7]\ _03903_ VPWR VGND _06889_ sg13g2_nor2_1
X_26626_ _03816_ _12524_ VPWR VGND _06890_ sg13g2_nor2_1
X_26627_ _12549_ _03819_ VPWR VGND _06891_ sg13g2_nor2_1
X_26628_ _04035_ _06890_ _06891_ _03911_ VPWR VGND 
+ _06892_
+ sg13g2_a22oi_1
X_26629_ _12524_ _03916_ VPWR VGND _06893_ sg13g2_nand2b_1
X_26630_ _03930_ _12549_ _06893_ VPWR VGND _06894_ sg13g2_o21ai_1
X_26631_ _03825_ _06894_ _04142_ VPWR VGND _06895_ sg13g2_a21oi_1
X_26632_ _03812_ _06892_ _06895_ VPWR VGND _06896_ sg13g2_a21oi_1
X_26633_ _04074_ _06888_ _06889_ _06896_ VPWR VGND 
+ _06897_
+ sg13g2_nor4_1
X_26634_ \atbs_core_0.spike_memory_0.n2417_o[7]\ _03804_ VPWR VGND _06898_ sg13g2_nor2_1
X_26635_ \atbs_core_0.spike_memory_0.n2414_o[7]\ _04702_ _03966_ VPWR VGND _06899_ sg13g2_o21ai_1
X_26636_ _04283_ _12581_ VPWR VGND _06900_ sg13g2_nor2_1
X_26637_ _12603_ _03852_ VPWR VGND _06901_ sg13g2_nor2_1
X_26638_ _04381_ _06900_ _06901_ _04343_ VPWR VGND 
+ _06902_
+ sg13g2_a22oi_1
X_26639_ _12581_ _04589_ VPWR VGND _06903_ sg13g2_nand2b_1
X_26640_ _04708_ _12603_ _06903_ VPWR VGND _06904_ sg13g2_o21ai_1
X_26641_ _03861_ _06904_ _03869_ VPWR VGND _06905_ sg13g2_a21oi_1
X_26642_ _04393_ _06902_ _06905_ VPWR VGND _06906_ sg13g2_a21oi_1
X_26643_ _06898_ _06899_ _06906_ VPWR VGND _06907_ sg13g2_nor3_1
X_26644_ \atbs_core_0.spike_memory_0.n2436_q[1204]\ _03804_ VPWR VGND _06908_ sg13g2_nor2_1
X_26645_ \atbs_core_0.spike_memory_0.n2418_o[7]\ _03946_ VPWR VGND _06909_ sg13g2_nor2_1
X_26646_ _03848_ _12637_ VPWR VGND _06910_ sg13g2_nor2_1
X_26647_ _12662_ _03852_ VPWR VGND _06911_ sg13g2_nor2_1
X_26648_ _03844_ _06910_ _06911_ _03857_ VPWR VGND 
+ _06912_
+ sg13g2_a22oi_1
X_26649_ _12637_ _03864_ VPWR VGND _06913_ sg13g2_nand2b_1
X_26650_ _04598_ _12662_ _06913_ VPWR VGND _06914_ sg13g2_o21ai_1
X_26651_ _03956_ _06914_ _04317_ VPWR VGND _06915_ sg13g2_a21oi_1
X_26652_ _03841_ _06912_ _06915_ VPWR VGND _06916_ sg13g2_a21oi_1
X_26653_ _12095_ _06908_ _06909_ _06916_ VPWR VGND 
+ _06917_
+ sg13g2_nor4_1
X_26654_ _06897_ _06907_ _06917_ VPWR VGND _06918_ sg13g2_nor3_1
X_26655_ \atbs_core_0.spike_memory_0.n2385_o[7]\ _03970_ VPWR VGND _06919_ sg13g2_nand2b_1
X_26656_ \atbs_core_0.spike_memory_0.n2382_o[7]\ _04771_ _06919_ VPWR VGND _06920_ sg13g2_o21ai_1
X_26657_ _03746_ _02295_ VPWR VGND _06921_ sg13g2_nor2_1
X_26658_ _02318_ _04006_ VPWR VGND _06922_ sg13g2_nor2_1
X_26659_ _03743_ _06921_ _06922_ _04512_ VPWR VGND 
+ _06923_
+ sg13g2_a22oi_1
X_26660_ _02295_ _04110_ VPWR VGND _06924_ sg13g2_nand2b_1
X_26661_ _04237_ _02318_ _06924_ VPWR VGND _06925_ sg13g2_o21ai_1
X_26662_ _04386_ _06925_ _04391_ VPWR VGND _06926_ sg13g2_a21oi_1
X_26663_ _04324_ _06923_ _06926_ VPWR VGND _06927_ sg13g2_a21oi_1
X_26664_ _06920_ _06927_ VPWR VGND _06928_ sg13g2_or2_1
X_26665_ \atbs_core_0.spike_memory_0.n2381_o[7]\ _12085_ VPWR VGND _06929_ sg13g2_nor2_1
X_26666_ \atbs_core_0.spike_memory_0.n2378_o[7]\ _04292_ VPWR VGND _06930_ sg13g2_nor2_1
X_26667_ _03854_ _02240_ VPWR VGND _06931_ sg13g2_nor2_1
X_26668_ _02263_ _03784_ VPWR VGND _06932_ sg13g2_nor2_1
X_26669_ _05245_ _06931_ _06932_ _03815_ VPWR VGND 
+ _06933_
+ sg13g2_a22oi_1
X_26670_ _02240_ _04455_ VPWR VGND _06934_ sg13g2_nand2b_1
X_26671_ _04050_ _02263_ _06934_ VPWR VGND _06935_ sg13g2_o21ai_1
X_26672_ _03757_ _06935_ _03867_ VPWR VGND _06936_ sg13g2_a21oi_1
X_26673_ _03992_ _06933_ _06936_ VPWR VGND _06937_ sg13g2_a21oi_1
X_26674_ _03726_ _06929_ _06930_ _06937_ VPWR VGND 
+ _06938_
+ sg13g2_nor4_1
X_26675_ \atbs_core_0.spike_memory_0.n2389_o[7]\ _03802_ VPWR VGND _06939_ sg13g2_nor2_1
X_26676_ \atbs_core_0.spike_memory_0.n2386_o[7]\ _04078_ VPWR VGND _06940_ sg13g2_nor2_1
X_26677_ _03988_ _02349_ VPWR VGND _06941_ sg13g2_nor2_1
X_26678_ _02373_ _03850_ VPWR VGND _06942_ sg13g2_nor2_1
X_26679_ _04062_ _06941_ _06942_ _04597_ VPWR VGND 
+ _06943_
+ sg13g2_a22oi_1
X_26680_ _02349_ _03981_ VPWR VGND _06944_ sg13g2_nand2b_1
X_26681_ _03846_ _02373_ _06944_ VPWR VGND _06945_ sg13g2_o21ai_1
X_26682_ _03859_ _06945_ _04068_ VPWR VGND _06946_ sg13g2_a21oi_1
X_26683_ _03839_ _06943_ _06946_ VPWR VGND _06947_ sg13g2_a21oi_1
X_26684_ _04746_ _06939_ _06940_ _06947_ VPWR VGND 
+ _06948_
+ sg13g2_nor4_1
X_26685_ _06938_ _06948_ _04276_ VPWR VGND _06949_ sg13g2_o21ai_1
X_26686_ _03924_ _06928_ _06949_ VPWR VGND _06950_ sg13g2_o21ai_1
X_26687_ \atbs_core_0.spike_memory_0.n2405_o[7]\ _04759_ VPWR VGND _06951_ sg13g2_nor2_1
X_26688_ \atbs_core_0.spike_memory_0.n2402_o[7]\ _03779_ VPWR VGND _06952_ sg13g2_nor2_1
X_26689_ _04254_ _02578_ VPWR VGND _06953_ sg13g2_nor2_1
X_26690_ _02599_ _03842_ VPWR VGND _06954_ sg13g2_nor2_1
X_26691_ _04108_ _06953_ _06954_ _03983_ VPWR VGND 
+ _06955_
+ sg13g2_a22oi_1
X_26692_ _02578_ _03988_ VPWR VGND _06956_ sg13g2_nand2b_1
X_26693_ _04425_ _02599_ _06956_ VPWR VGND _06957_ sg13g2_o21ai_1
X_26694_ _05510_ _06957_ _03810_ VPWR VGND _06958_ sg13g2_a21oi_1
X_26695_ _04118_ _06955_ _06958_ VPWR VGND _06959_ sg13g2_a21oi_1
X_26696_ _12093_ _06951_ _06952_ _06959_ VPWR VGND 
+ _06960_
+ sg13g2_nor4_1
X_26697_ \atbs_core_0.spike_memory_0.n2401_o[7]\ _12086_ VPWR VGND _06961_ sg13g2_nor2_1
X_26698_ \atbs_core_0.spike_memory_0.n2398_o[7]\ _04000_ _03722_ VPWR VGND _06962_ sg13g2_o21ai_1
X_26699_ _03787_ _02531_ VPWR VGND _06963_ sg13g2_nor2_1
X_26700_ _02552_ _03785_ VPWR VGND _06964_ sg13g2_nor2_1
X_26701_ _03782_ _06963_ _06964_ _03754_ VPWR VGND 
+ _06965_
+ sg13g2_a22oi_1
X_26702_ _02531_ _03891_ VPWR VGND _06966_ sg13g2_nand2b_1
X_26703_ _03753_ _02552_ _06966_ VPWR VGND _06967_ sg13g2_o21ai_1
X_26704_ _03758_ _06967_ _04294_ VPWR VGND _06968_ sg13g2_a21oi_1
X_26705_ _03739_ _06965_ _06968_ VPWR VGND _06969_ sg13g2_a21oi_1
X_26706_ _06961_ _06962_ _06969_ VPWR VGND _06970_ sg13g2_nor3_1
X_26707_ \atbs_core_0.spike_memory_0.n2397_o[7]\ _04759_ VPWR VGND _06971_ sg13g2_nor2_1
X_26708_ \atbs_core_0.spike_memory_0.n2394_o[7]\ _03779_ VPWR VGND _06972_ sg13g2_nor2_1
X_26709_ _04237_ _02482_ VPWR VGND _06973_ sg13g2_nor2_1
X_26710_ _02504_ _04006_ VPWR VGND _06974_ sg13g2_nor2_1
X_26711_ _04003_ _06973_ _06974_ _03978_ VPWR VGND 
+ _06975_
+ sg13g2_a22oi_1
X_26712_ _02482_ _04110_ VPWR VGND _06976_ sg13g2_nand2b_1
X_26713_ _04004_ _02504_ _06976_ VPWR VGND _06977_ sg13g2_o21ai_1
X_26714_ _04386_ _06977_ _03839_ VPWR VGND _06978_ sg13g2_a21oi_1
X_26715_ _04324_ _06975_ _06978_ VPWR VGND _06979_ sg13g2_a21oi_1
X_26716_ _03727_ _06971_ _06972_ _06979_ VPWR VGND 
+ _06980_
+ sg13g2_nor4_1
X_26717_ _06960_ _06970_ _06980_ VPWR VGND _06981_ sg13g2_or3_1
X_26718_ _03720_ _06950_ _06981_ _03717_ _04335_ VPWR 
+ VGND
+ _06982_ sg13g2_a221oi_1
X_26719_ _12079_ _06918_ _06982_ VPWR VGND _06983_ sg13g2_o21ai_1
X_26720_ _04503_ _06887_ _06983_ VPWR VGND _06984_ sg13g2_nand3_1
X_26721_ _04333_ _06860_ _06984_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[7]\ sg13g2_o21ai_1
X_26722_ _03747_ _02399_ VPWR VGND _06985_ sg13g2_nor2_1
X_26723_ _02418_ _03751_ VPWR VGND _06986_ sg13g2_nor2_1
X_26724_ _03744_ _06985_ _06986_ _03755_ VPWR VGND 
+ _06987_
+ sg13g2_a22oi_1
X_26725_ _02399_ _03764_ VPWR VGND _06988_ sg13g2_nand2b_1
X_26726_ _03761_ _02418_ _06988_ VPWR VGND _06989_ sg13g2_o21ai_1
X_26727_ _03759_ _06989_ _03769_ VPWR VGND _06990_ sg13g2_a21oi_1
X_26728_ _03740_ _06987_ _06990_ VPWR VGND _06991_ sg13g2_a21oi_1
X_26729_ _00135_ _03733_ _03737_ _02448_ _06991_ VPWR 
+ VGND
+ _06992_ sg13g2_a221oi_1
X_26730_ \atbs_core_0.spike_memory_0.n2401_o[8]\ _03776_ VPWR VGND _06993_ sg13g2_nor2_1
X_26731_ \atbs_core_0.spike_memory_0.n2398_o[8]\ _03779_ _03780_ VPWR VGND _06994_ sg13g2_o21ai_1
X_26732_ _02711_ _02532_ VPWR VGND _06995_ sg13g2_nor2_1
X_26733_ _02553_ _03785_ VPWR VGND _06996_ sg13g2_nor2_1
X_26734_ _03782_ _06995_ _06996_ _03788_ VPWR VGND 
+ _06997_
+ sg13g2_a22oi_1
X_26735_ _02532_ _03891_ VPWR VGND _06998_ sg13g2_nand2b_1
X_26736_ _03746_ _02553_ _06998_ VPWR VGND _06999_ sg13g2_o21ai_1
X_26737_ _03790_ _06999_ _03768_ VPWR VGND _07000_ sg13g2_a21oi_1
X_26738_ _02700_ _06997_ _07000_ VPWR VGND _07001_ sg13g2_a21oi_1
X_26739_ _06993_ _06994_ _07001_ VPWR VGND _07002_ sg13g2_or3_1
X_26740_ _03775_ _07002_ VPWR VGND _07003_ sg13g2_nand2_1
X_26741_ _03729_ _06992_ _07003_ VPWR VGND _07004_ sg13g2_o21ai_1
X_26742_ \atbs_core_0.spike_memory_0.n2397_o[8]\ _03804_ VPWR VGND _07005_ sg13g2_nor2_1
X_26743_ \atbs_core_0.spike_memory_0.n2394_o[8]\ _03807_ VPWR VGND _07006_ sg13g2_nor2_1
X_26744_ _03816_ _02485_ VPWR VGND _07007_ sg13g2_nor2_1
X_26745_ _02506_ _03819_ VPWR VGND _07008_ sg13g2_nor2_1
X_26746_ _04035_ _07007_ _07008_ _03823_ VPWR VGND 
+ _07009_
+ sg13g2_a22oi_1
X_26747_ _02485_ _03916_ VPWR VGND _07010_ sg13g2_nand2b_1
X_26748_ _03826_ _02506_ _07010_ VPWR VGND _07011_ sg13g2_o21ai_1
X_26749_ _03825_ _07011_ _03831_ VPWR VGND _07012_ sg13g2_a21oi_1
X_26750_ _03812_ _07009_ _07012_ VPWR VGND _07013_ sg13g2_a21oi_1
X_26751_ _07005_ _07006_ _07013_ VPWR VGND _07014_ sg13g2_nor3_1
X_26752_ \atbs_core_0.spike_memory_0.n2405_o[8]\ _03736_ VPWR VGND _07015_ sg13g2_nand2b_1
X_26753_ \atbs_core_0.spike_memory_0.n2402_o[8]\ _03836_ _07015_ VPWR VGND _07016_ sg13g2_o21ai_1
X_26754_ _03848_ _02579_ VPWR VGND _07017_ sg13g2_nor2_1
X_26755_ _02600_ _03852_ VPWR VGND _07018_ sg13g2_nor2_1
X_26756_ _03844_ _07017_ _07018_ _03857_ VPWR VGND 
+ _07019_
+ sg13g2_a22oi_1
X_26757_ _02579_ _03864_ VPWR VGND _07020_ sg13g2_nand2b_1
X_26758_ _03856_ _02600_ _07020_ VPWR VGND _07021_ sg13g2_o21ai_1
X_26759_ _03861_ _07021_ _03869_ VPWR VGND _07022_ sg13g2_a21oi_1
X_26760_ _03841_ _07019_ _07022_ VPWR VGND _07023_ sg13g2_a21oi_1
X_26761_ _07016_ _07023_ _03872_ VPWR VGND _07024_ sg13g2_o21ai_1
X_26762_ _03801_ _07014_ _07024_ VPWR VGND _07025_ sg13g2_o21ai_1
X_26763_ _03725_ _07004_ _07025_ _07002_ VPWR VGND 
+ _07026_
+ sg13g2_a22oi_1
X_26764_ \atbs_core_0.spike_memory_0.n2365_o[8]\ _03877_ VPWR VGND _07027_ sg13g2_nor2_1
X_26765_ \atbs_core_0.spike_memory_0.n2362_o[8]\ _03836_ VPWR VGND _07028_ sg13g2_nor2_1
X_26766_ _03882_ _12556_ VPWR VGND _07029_ sg13g2_nor2_1
X_26767_ _02008_ _04023_ VPWR VGND _07030_ sg13g2_nor2_1
X_26768_ _03881_ _07029_ _07030_ _03887_ VPWR VGND 
+ _07031_
+ sg13g2_a22oi_1
X_26769_ _12556_ _04026_ VPWR VGND _07032_ sg13g2_nand2b_1
X_26770_ _03886_ _02008_ _07032_ VPWR VGND _07033_ sg13g2_o21ai_1
X_26771_ _03889_ _07033_ _03895_ VPWR VGND _07034_ sg13g2_a21oi_1
X_26772_ _03880_ _07031_ _07034_ VPWR VGND _07035_ sg13g2_a21oi_1
X_26773_ _03728_ _07027_ _07028_ _07035_ VPWR VGND 
+ _07036_
+ sg13g2_nor4_1
X_26774_ \atbs_core_0.spike_memory_0.n2373_o[8]\ _12087_ VPWR VGND _07037_ sg13g2_nor2_1
X_26775_ \atbs_core_0.spike_memory_0.n2370_o[8]\ _03903_ VPWR VGND _07038_ sg13g2_nor2_1
X_26776_ _03907_ _02089_ VPWR VGND _07039_ sg13g2_nor2_1
X_26777_ _02112_ _03909_ VPWR VGND _07040_ sg13g2_nor2_1
X_26778_ _03906_ _07039_ _07040_ _03911_ VPWR VGND 
+ _07041_
+ sg13g2_a22oi_1
X_26779_ _02089_ _05745_ VPWR VGND _07042_ sg13g2_nand2b_1
X_26780_ _03914_ _02112_ _07042_ VPWR VGND _07043_ sg13g2_o21ai_1
X_26781_ _03913_ _07043_ _03919_ VPWR VGND _07044_ sg13g2_a21oi_1
X_26782_ _03905_ _07041_ _07044_ VPWR VGND _07045_ sg13g2_a21oi_1
X_26783_ _03900_ _07037_ _07038_ _07045_ VPWR VGND 
+ _07046_
+ sg13g2_nor4_1
X_26784_ _03724_ _07036_ _07046_ VPWR VGND _07047_ sg13g2_nor3_1
X_26785_ \atbs_core_0.spike_memory_0.n2361_o[8]\ _12087_ VPWR VGND _07048_ sg13g2_nor2_1
X_26786_ \atbs_core_0.spike_memory_0.n2358_o[8]\ _04702_ VPWR VGND _07049_ sg13g2_nor2_1
X_26787_ _03930_ _02118_ VPWR VGND _07050_ sg13g2_nor2_1
X_26788_ _02285_ _03932_ VPWR VGND _07051_ sg13g2_nor2_1
X_26789_ _03929_ _07050_ _07051_ _02713_ VPWR VGND 
+ _07052_
+ sg13g2_a22oi_1
X_26790_ _02118_ _03937_ VPWR VGND _07053_ sg13g2_nand2b_1
X_26791_ _02712_ _02285_ _07053_ VPWR VGND _07054_ sg13g2_o21ai_1
X_26792_ _03889_ _07054_ _04263_ VPWR VGND _07055_ sg13g2_a21oi_1
X_26793_ _02701_ _07052_ _07055_ VPWR VGND _07056_ sg13g2_a21oi_1
X_26794_ _03728_ _07048_ _07049_ _07056_ VPWR VGND 
+ _07057_
+ sg13g2_nor4_1
X_26795_ \atbs_core_0.spike_memory_0.n2369_o[8]\ _03901_ VPWR VGND _07058_ sg13g2_nor2_1
X_26796_ \atbs_core_0.spike_memory_0.n2366_o[8]\ _03807_ VPWR VGND _07059_ sg13g2_nor2_1
X_26797_ _04052_ _02034_ VPWR VGND _07060_ sg13g2_nor2_1
X_26798_ _02055_ _03952_ VPWR VGND _07061_ sg13g2_nor2_1
X_26799_ _03814_ _07060_ _07061_ _03823_ VPWR VGND 
+ _07062_
+ sg13g2_a22oi_1
X_26800_ _02034_ _03827_ VPWR VGND _07063_ sg13g2_nand2b_1
X_26801_ _03816_ _02055_ _07063_ VPWR VGND _07064_ sg13g2_o21ai_1
X_26802_ _03825_ _07064_ _03831_ VPWR VGND _07065_ sg13g2_a21oi_1
X_26803_ _03948_ _07062_ _07065_ VPWR VGND _07066_ sg13g2_a21oi_1
X_26804_ _03900_ _07058_ _07059_ _07066_ VPWR VGND 
+ _07067_
+ sg13g2_nor4_1
X_26805_ _03925_ _07057_ _07067_ VPWR VGND _07068_ sg13g2_nor3_1
X_26806_ _07047_ _07068_ _03721_ VPWR VGND _07069_ sg13g2_o21ai_1
X_26807_ _03721_ _07026_ _07069_ VPWR VGND _07070_ sg13g2_o21ai_1
X_26808_ _03821_ _02144_ VPWR VGND _07071_ sg13g2_nor2_1
X_26809_ _02167_ _03818_ VPWR VGND _07072_ sg13g2_nor2_1
X_26810_ _03813_ _07071_ _07072_ _03914_ VPWR VGND 
+ _07073_
+ sg13g2_a22oi_1
X_26811_ _02144_ _03791_ VPWR VGND _07074_ sg13g2_nand2b_1
X_26812_ _02711_ _02167_ _07074_ VPWR VGND _07075_ sg13g2_o21ai_1
X_26813_ _03790_ _07075_ _03830_ VPWR VGND _07076_ sg13g2_a21oi_1
X_26814_ _02700_ _07073_ _07076_ VPWR VGND _07077_ sg13g2_a21oi_1
X_26815_ _00136_ _03732_ _03736_ _02200_ _07077_ VPWR 
+ VGND
+ _07078_ sg13g2_a221oi_1
X_26816_ \atbs_core_0.spike_memory_0.n2385_o[8]\ _03802_ VPWR VGND _07079_ sg13g2_nor2_1
X_26817_ \atbs_core_0.spike_memory_0.n2382_o[8]\ _03778_ _07552_ VPWR VGND _07080_ sg13g2_o21ai_1
X_26818_ _04050_ _02296_ VPWR VGND _07081_ sg13g2_nor2_1
X_26819_ _02319_ _03784_ VPWR VGND _07082_ sg13g2_nor2_1
X_26820_ _05245_ _07081_ _07082_ _03821_ VPWR VGND 
+ _07083_
+ sg13g2_a22oi_1
X_26821_ _02296_ _04455_ VPWR VGND _07084_ sg13g2_nand2b_1
X_26822_ _03745_ _02319_ _07084_ VPWR VGND _07085_ sg13g2_o21ai_1
X_26823_ _03757_ _07085_ _03867_ VPWR VGND _07086_ sg13g2_a21oi_1
X_26824_ _03810_ _07083_ _07086_ VPWR VGND _07087_ sg13g2_a21oi_1
X_26825_ _07079_ _07080_ _07087_ VPWR VGND _07088_ sg13g2_or3_1
X_26826_ _03774_ _07088_ VPWR VGND _07089_ sg13g2_nand2_1
X_26827_ _03926_ _07078_ _07089_ VPWR VGND _07090_ sg13g2_o21ai_1
X_26828_ \atbs_core_0.spike_memory_0.n2381_o[8]\ _04245_ VPWR VGND _07091_ sg13g2_nor2_1
X_26829_ \atbs_core_0.spike_memory_0.n2378_o[8]\ _04247_ VPWR VGND _07092_ sg13g2_nor2_1
X_26830_ _05533_ _02241_ VPWR VGND _07093_ sg13g2_nor2_1
X_26831_ _02264_ _03851_ VPWR VGND _07094_ sg13g2_nor2_1
X_26832_ _03843_ _07093_ _07094_ _04708_ VPWR VGND 
+ _07095_
+ sg13g2_a22oi_1
X_26833_ _02241_ _03982_ VPWR VGND _07096_ sg13g2_nand2b_1
X_26834_ _03847_ _02264_ _07096_ VPWR VGND _07097_ sg13g2_o21ai_1
X_26835_ _03860_ _07097_ _04287_ VPWR VGND _07098_ sg13g2_a21oi_1
X_26836_ _03840_ _07095_ _07098_ VPWR VGND _07099_ sg13g2_a21oi_1
X_26837_ _07091_ _07092_ _07099_ VPWR VGND _07100_ sg13g2_nor3_1
X_26838_ \atbs_core_0.spike_memory_0.n2389_o[8]\ _03735_ VPWR VGND _07101_ sg13g2_nand2b_1
X_26839_ \atbs_core_0.spike_memory_0.n2386_o[8]\ _05540_ _07101_ VPWR VGND _07102_ sg13g2_o21ai_1
X_26840_ _04267_ _02350_ VPWR VGND _07103_ sg13g2_nor2_1
X_26841_ _02375_ _04250_ VPWR VGND _07104_ sg13g2_nor2_1
X_26842_ _04023_ _07103_ _07104_ _04090_ VPWR VGND 
+ _07105_
+ sg13g2_a22oi_1
X_26843_ _02350_ _03977_ VPWR VGND _07106_ sg13g2_nand2b_1
X_26844_ _04089_ _02375_ _07106_ VPWR VGND _07107_ sg13g2_o21ai_1
X_26845_ _04253_ _07107_ _04272_ VPWR VGND _07108_ sg13g2_a21oi_1
X_26846_ _03895_ _07105_ _07108_ VPWR VGND _07109_ sg13g2_a21oi_1
X_26847_ _07102_ _07109_ _03774_ VPWR VGND _07110_ sg13g2_o21ai_1
X_26848_ _04074_ _07100_ _07110_ VPWR VGND _07111_ sg13g2_o21ai_1
X_26849_ _03724_ _07090_ _07111_ _07088_ VPWR VGND 
+ _07112_
+ sg13g2_a22oi_1
X_26850_ _04045_ _07112_ VPWR VGND _07113_ sg13g2_and2_1
X_26851_ _03761_ _02627_ VPWR VGND _07114_ sg13g2_nor2_1
X_26852_ _02648_ _04280_ VPWR VGND _07115_ sg13g2_nor2_1
X_26853_ _04510_ _07114_ _07115_ _04513_ VPWR VGND 
+ _07116_
+ sg13g2_a22oi_1
X_26854_ _02627_ _04267_ VPWR VGND _07117_ sg13g2_nand2b_1
X_26855_ _03978_ _02648_ _07117_ VPWR VGND _07118_ sg13g2_o21ai_1
X_26856_ _04387_ _07118_ _03840_ VPWR VGND _07119_ sg13g2_a21oi_1
X_26857_ _04376_ _07116_ _07119_ VPWR VGND _07120_ sg13g2_a21oi_1
X_26858_ _00134_ _03969_ _03972_ _02676_ _07120_ VPWR 
+ VGND
+ _07121_ sg13g2_a221oi_1
X_26859_ \atbs_core_0.spike_memory_0.n2417_o[8]\ _12086_ VPWR VGND _07122_ sg13g2_nor2_1
X_26860_ \atbs_core_0.spike_memory_0.n2414_o[8]\ _04771_ _03722_ VPWR VGND _07123_ sg13g2_o21ai_1
X_26861_ _03746_ _12582_ VPWR VGND _07124_ sg13g2_nor2_1
X_26862_ _12605_ _03750_ VPWR VGND _07125_ sg13g2_nor2_1
X_26863_ _03743_ _07124_ _07125_ _03761_ VPWR VGND 
+ _07126_
+ sg13g2_a22oi_1
X_26864_ _12582_ _03763_ VPWR VGND _07127_ sg13g2_nand2b_1
X_26865_ _04115_ _12605_ _07127_ VPWR VGND _07128_ sg13g2_o21ai_1
X_26866_ _03758_ _07128_ _04294_ VPWR VGND _07129_ sg13g2_a21oi_1
X_26867_ _03739_ _07126_ _07129_ VPWR VGND _07130_ sg13g2_a21oi_1
X_26868_ _07122_ _07123_ _07130_ VPWR VGND _07131_ sg13g2_or3_1
X_26869_ _03775_ _07131_ VPWR VGND _07132_ sg13g2_nand2_1
X_26870_ _03729_ _07121_ _07132_ VPWR VGND _07133_ sg13g2_o21ai_1
X_26871_ \atbs_core_0.spike_memory_0.n2413_o[8]\ _03944_ VPWR VGND _07134_ sg13g2_nor2_1
X_26872_ \atbs_core_0.spike_memory_0.n2410_o[8]\ _03807_ VPWR VGND _07135_ sg13g2_nor2_1
X_26873_ _03822_ _12527_ VPWR VGND _07136_ sg13g2_nor2_1
X_26874_ _12550_ _03909_ VPWR VGND _07137_ sg13g2_nor2_1
X_26875_ _04150_ _07136_ _07137_ _04154_ VPWR VGND 
+ _07138_
+ sg13g2_a22oi_1
X_26876_ _12527_ _05745_ VPWR VGND _07139_ sg13g2_nand2b_1
X_26877_ _05753_ _12550_ _07139_ VPWR VGND _07140_ sg13g2_o21ai_1
X_26878_ _03913_ _07140_ _03919_ VPWR VGND _07141_ sg13g2_a21oi_1
X_26879_ _03905_ _07138_ _07141_ VPWR VGND _07142_ sg13g2_a21oi_1
X_26880_ _07134_ _07135_ _07142_ VPWR VGND _07143_ sg13g2_nor3_1
X_26881_ \atbs_core_0.spike_memory_0.n2436_q[1205]\ _03971_ VPWR VGND _07144_ sg13g2_nand2b_1
X_26882_ \atbs_core_0.spike_memory_0.n2418_o[8]\ _04527_ _07144_ VPWR VGND _07145_ sg13g2_o21ai_1
X_26883_ _03856_ _12638_ VPWR VGND _07146_ sg13g2_nor2_1
X_26884_ _12663_ _03952_ VPWR VGND _07147_ sg13g2_nor2_1
X_26885_ _03844_ _07146_ _07147_ _03823_ VPWR VGND 
+ _07148_
+ sg13g2_a22oi_1
X_26886_ _12638_ _04167_ VPWR VGND _07149_ sg13g2_nand2b_1
X_26887_ _03949_ _12663_ _07149_ VPWR VGND _07150_ sg13g2_o21ai_1
X_26888_ _03956_ _07150_ _04317_ VPWR VGND _07151_ sg13g2_a21oi_1
X_26889_ _03948_ _07148_ _07151_ VPWR VGND _07152_ sg13g2_a21oi_1
X_26890_ _07145_ _07152_ _03775_ VPWR VGND _07153_ sg13g2_o21ai_1
X_26891_ _03801_ _07143_ _07153_ VPWR VGND _07154_ sg13g2_o21ai_1
X_26892_ _03725_ _07133_ _07154_ _07131_ _03721_ VPWR 
+ VGND
+ _07155_ sg13g2_a221oi_1
X_26893_ _03718_ _07113_ _07155_ VPWR VGND _07156_ sg13g2_nor3_1
X_26894_ _03719_ _07070_ _07156_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[8]\ sg13g2_a21oi_1
X_26895_ _04340_ _02400_ VPWR VGND _07157_ sg13g2_nor2_1
X_26896_ _02419_ _03976_ VPWR VGND _07158_ sg13g2_nor2_1
X_26897_ _04339_ _07157_ _07158_ _04343_ VPWR VGND 
+ _07159_
+ sg13g2_a22oi_1
X_26898_ _02400_ _03788_ VPWR VGND _07160_ sg13g2_nand2b_1
X_26899_ _04347_ _02419_ _07160_ VPWR VGND _07161_ sg13g2_o21ai_1
X_26900_ _04345_ _07161_ _03974_ VPWR VGND _07162_ sg13g2_a21oi_1
X_26901_ _04338_ _07159_ _07162_ VPWR VGND _07163_ sg13g2_a21oi_1
X_26902_ _00138_ _03733_ _03737_ _02450_ _07163_ VPWR 
+ VGND
+ _07164_ sg13g2_a221oi_1
X_26903_ _04357_ _02145_ VPWR VGND _07165_ sg13g2_nor2_1
X_26904_ _02168_ _04359_ VPWR VGND _07166_ sg13g2_nor2_1
X_26905_ _04356_ _07165_ _07166_ _04362_ VPWR VGND 
+ _07167_
+ sg13g2_a22oi_1
X_26906_ _02145_ _03907_ VPWR VGND _07168_ sg13g2_nand2b_1
X_26907_ _04365_ _02168_ _07168_ VPWR VGND _07169_ sg13g2_o21ai_1
X_26908_ _04364_ _07169_ _04021_ VPWR VGND _07170_ sg13g2_a21oi_1
X_26909_ _04355_ _07167_ _07170_ VPWR VGND _07171_ sg13g2_a21oi_1
X_26910_ _00139_ _04353_ _04354_ _02205_ _07171_ VPWR 
+ VGND
+ _07172_ sg13g2_a221oi_1
X_26911_ _04337_ _07164_ _07172_ _04371_ _04688_ VPWR 
+ VGND
+ _07173_ sg13g2_a221oi_1
X_26912_ _02713_ _02628_ VPWR VGND _07174_ sg13g2_nor2_1
X_26913_ _02649_ _04533_ VPWR VGND _07175_ sg13g2_nor2_1
X_26914_ _04531_ _07174_ _07175_ _04536_ VPWR VGND 
+ _07176_
+ sg13g2_a22oi_1
X_26915_ _02628_ _04320_ VPWR VGND _07177_ sg13g2_nand2b_1
X_26916_ _03887_ _02649_ _07177_ VPWR VGND _07178_ sg13g2_o21ai_1
X_26917_ _04538_ _07178_ _04542_ VPWR VGND _07179_ sg13g2_a21oi_1
X_26918_ _04530_ _07176_ _07179_ VPWR VGND _07180_ sg13g2_a21oi_1
X_26919_ _00137_ _04660_ _04661_ _02678_ _07180_ VPWR 
+ VGND
+ _07181_ sg13g2_a221oi_1
X_26920_ _05483_ _07181_ VPWR VGND _07182_ sg13g2_nand2_1
X_26921_ \atbs_core_0.spike_memory_0.n2385_o[9]\ _03735_ VPWR VGND _07183_ sg13g2_nand2b_1
X_26922_ \atbs_core_0.spike_memory_0.n2382_o[9]\ _04102_ _07183_ VPWR VGND _07184_ sg13g2_o21ai_1
X_26923_ _04346_ _02297_ VPWR VGND _07185_ sg13g2_nor2_1
X_26924_ _02320_ _04265_ VPWR VGND _07186_ sg13g2_nor2_1
X_26925_ _05496_ _07185_ _07186_ _04268_ VPWR VGND 
+ _07187_
+ sg13g2_a22oi_1
X_26926_ _02297_ _03760_ VPWR VGND _07188_ sg13g2_nand2b_1
X_26927_ _04267_ _02320_ _07188_ VPWR VGND _07189_ sg13g2_o21ai_1
X_26928_ _04235_ _07189_ _03973_ VPWR VGND _07190_ sg13g2_a21oi_1
X_26929_ _03940_ _07187_ _07190_ VPWR VGND _07191_ sg13g2_a21oi_1
X_26930_ _07184_ _07191_ VPWR VGND _07192_ sg13g2_or2_1
X_26931_ \atbs_core_0.spike_memory_0.n2381_o[9]\ _04075_ VPWR VGND _07193_ sg13g2_nor2_1
X_26932_ \atbs_core_0.spike_memory_0.n2378_o[9]\ _04229_ VPWR VGND _07194_ sg13g2_nor2_1
X_26933_ _04054_ _02242_ VPWR VGND _07195_ sg13g2_nor2_1
X_26934_ _02265_ _03742_ VPWR VGND _07196_ sg13g2_nor2_1
X_26935_ _04422_ _07195_ _07196_ _03827_ VPWR VGND 
+ _07197_
+ sg13g2_a22oi_1
X_26936_ _02242_ _03745_ VPWR VGND _07198_ sg13g2_nand2b_1
X_26937_ _03915_ _02265_ _07198_ VPWR VGND _07199_ sg13g2_o21ai_1
X_26938_ _03986_ _07199_ _03738_ VPWR VGND _07200_ sg13g2_a21oi_1
X_26939_ _04839_ _07197_ _07200_ VPWR VGND _07201_ sg13g2_a21oi_1
X_26940_ _03773_ _07193_ _07194_ _07201_ VPWR VGND 
+ _07202_
+ sg13g2_nor4_1
X_26941_ \atbs_core_0.spike_memory_0.n2389_o[9]\ _04075_ VPWR VGND _07203_ sg13g2_nor2_1
X_26942_ \atbs_core_0.spike_memory_0.n2386_o[9]\ _04000_ VPWR VGND _07204_ sg13g2_nor2_1
X_26943_ _03863_ _02353_ VPWR VGND _07205_ sg13g2_nor2_1
X_26944_ _02376_ _05245_ VPWR VGND _07206_ sg13g2_nor2_1
X_26945_ _04086_ _07205_ _07206_ _04167_ VPWR VGND 
+ _07207_
+ sg13g2_a22oi_1
X_26946_ _02353_ _03854_ VPWR VGND _07208_ sg13g2_nand2b_1
X_26947_ _04480_ _02376_ _07208_ VPWR VGND _07209_ sg13g2_o21ai_1
X_26948_ _05510_ _07209_ _03738_ VPWR VGND _07210_ sg13g2_a21oi_1
X_26949_ _04098_ _07207_ _07210_ VPWR VGND _07211_ sg13g2_a21oi_1
X_26950_ _04746_ _07203_ _07204_ _07211_ VPWR VGND 
+ _07212_
+ sg13g2_nor4_1
X_26951_ _07202_ _07212_ _03924_ VPWR VGND _07213_ sg13g2_o21ai_1
X_26952_ _04277_ _07192_ _07213_ VPWR VGND _07214_ sg13g2_o21ai_1
X_26953_ \atbs_core_0.spike_memory_0.n2405_o[9]\ _04245_ VPWR VGND _07215_ sg13g2_nor2_1
X_26954_ \atbs_core_0.spike_memory_0.n2402_o[9]\ _04247_ VPWR VGND _07216_ sg13g2_nor2_1
X_26955_ _04413_ _02580_ VPWR VGND _07217_ sg13g2_nor2_1
X_26956_ _02602_ _04422_ VPWR VGND _07218_ sg13g2_nor2_1
X_26957_ _04280_ _07217_ _07218_ _04704_ VPWR VGND 
+ _07219_
+ sg13g2_a22oi_1
X_26958_ _02580_ _04425_ VPWR VGND _07220_ sg13g2_nand2b_1
X_26959_ _05533_ _02602_ _07220_ VPWR VGND _07221_ sg13g2_o21ai_1
X_26960_ _04092_ _07221_ _04287_ VPWR VGND _07222_ sg13g2_a21oi_1
X_26961_ _04392_ _07219_ _07222_ VPWR VGND _07223_ sg13g2_a21oi_1
X_26962_ _12094_ _07215_ _07216_ _07223_ VPWR VGND 
+ _07224_
+ sg13g2_nor4_1
X_26963_ \atbs_core_0.spike_memory_0.n2401_o[9]\ _04076_ VPWR VGND _07225_ sg13g2_nor2_1
X_26964_ \atbs_core_0.spike_memory_0.n2398_o[9]\ _05540_ _03723_ VPWR VGND _07226_ sg13g2_o21ai_1
X_26965_ _04026_ _02533_ VPWR VGND _07227_ sg13g2_nor2_1
X_26966_ _02554_ _04108_ VPWR VGND _07228_ sg13g2_nor2_1
X_26967_ _04152_ _07227_ _07228_ _05544_ VPWR VGND 
+ _07229_
+ sg13g2_a22oi_1
X_26968_ _02533_ _04115_ VPWR VGND _07230_ sg13g2_nand2b_1
X_26969_ _03764_ _02554_ _07230_ VPWR VGND _07231_ sg13g2_o21ai_1
X_26970_ _04114_ _07231_ _04118_ VPWR VGND _07232_ sg13g2_a21oi_1
X_26971_ _04142_ _07229_ _07232_ VPWR VGND _07233_ sg13g2_a21oi_1
X_26972_ _07225_ _07226_ _07233_ VPWR VGND _07234_ sg13g2_nor3_1
X_26973_ \atbs_core_0.spike_memory_0.n2397_o[9]\ _04260_ VPWR VGND _07235_ sg13g2_nor2_1
X_26974_ \atbs_core_0.spike_memory_0.n2394_o[9]\ _04079_ VPWR VGND _07236_ sg13g2_nor2_1
X_26975_ _04236_ _02486_ VPWR VGND _07237_ sg13g2_nor2_1
X_26976_ _02507_ _04250_ VPWR VGND _07238_ sg13g2_nor2_1
X_26977_ _03884_ _07237_ _07238_ _04518_ VPWR VGND 
+ _07239_
+ sg13g2_a22oi_1
X_26978_ _02486_ _04004_ VPWR VGND _07240_ sg13g2_nand2b_1
X_26979_ _04083_ _02507_ _07240_ VPWR VGND _07241_ sg13g2_o21ai_1
X_26980_ _04253_ _07241_ _04272_ VPWR VGND _07242_ sg13g2_a21oi_1
X_26981_ _03895_ _07239_ _07242_ VPWR VGND _07243_ sg13g2_a21oi_1
X_26982_ _04244_ _07235_ _07236_ _07243_ VPWR VGND 
+ _07244_
+ sg13g2_nor4_1
X_26983_ _07224_ _07234_ _07244_ VPWR VGND _07245_ sg13g2_or3_1
X_26984_ _04330_ _07214_ _07245_ _03718_ _04335_ VPWR 
+ VGND
+ _07246_ sg13g2_a221oi_1
X_26985_ \atbs_core_0.spike_memory_0.n2413_o[9]\ _04372_ VPWR VGND _07247_ sg13g2_nor2_1
X_26986_ \atbs_core_0.spike_memory_0.n2410_o[9]\ _04032_ VPWR VGND _07248_ sg13g2_nor2_1
X_26987_ _03747_ _12528_ VPWR VGND _07249_ sg13g2_nor2_1
X_26988_ _12551_ _03751_ VPWR VGND _07250_ sg13g2_nor2_1
X_26989_ _03744_ _07249_ _07250_ _04379_ VPWR VGND 
+ _07251_
+ sg13g2_a22oi_1
X_26990_ _12528_ _04111_ VPWR VGND _07252_ sg13g2_nand2b_1
X_26991_ _04512_ _12551_ _07252_ VPWR VGND _07253_ sg13g2_o21ai_1
X_26992_ _04387_ _07253_ _04392_ VPWR VGND _07254_ sg13g2_a21oi_1
X_26993_ _04376_ _07251_ _07254_ VPWR VGND _07255_ sg13g2_a21oi_1
X_26994_ _03800_ _07247_ _07248_ _07255_ VPWR VGND 
+ _07256_
+ sg13g2_nor4_1
X_26995_ \atbs_core_0.spike_memory_0.n2417_o[9]\ _03944_ VPWR VGND _07257_ sg13g2_nor2_1
X_26996_ \atbs_core_0.spike_memory_0.n2414_o[9]\ _04230_ _03723_ VPWR VGND _07258_ sg13g2_o21ai_1
X_26997_ _03822_ _12583_ VPWR VGND _07259_ sg13g2_nor2_1
X_26998_ _12606_ _03909_ VPWR VGND _07260_ sg13g2_nor2_1
X_26999_ _03906_ _07259_ _07260_ _04154_ VPWR VGND 
+ _07261_
+ sg13g2_a22oi_1
X_27000_ _12583_ _05745_ VPWR VGND _07262_ sg13g2_nand2b_1
X_27001_ _03914_ _12606_ _07262_ VPWR VGND _07263_ sg13g2_o21ai_1
X_27002_ _03913_ _07263_ _03919_ VPWR VGND _07264_ sg13g2_a21oi_1
X_27003_ _03905_ _07261_ _07264_ VPWR VGND _07265_ sg13g2_a21oi_1
X_27004_ _07257_ _07258_ _07265_ VPWR VGND _07266_ sg13g2_nor3_1
X_27005_ \atbs_core_0.spike_memory_0.n2436_q[1206]\ _03877_ VPWR VGND _07267_ sg13g2_nor2_1
X_27006_ \atbs_core_0.spike_memory_0.n2418_o[9]\ _04702_ VPWR VGND _07268_ sg13g2_nor2_1
X_27007_ _05753_ _12639_ VPWR VGND _07269_ sg13g2_nor2_1
X_27008_ _12665_ _05496_ VPWR VGND _07270_ sg13g2_nor2_1
X_27009_ _04628_ _07269_ _07270_ _04574_ VPWR VGND 
+ _07271_
+ sg13g2_a22oi_1
X_27010_ _12639_ _03892_ VPWR VGND _07272_ sg13g2_nand2b_1
X_27011_ _03882_ _12665_ _07272_ VPWR VGND _07273_ sg13g2_o21ai_1
X_27012_ _03889_ _07273_ _04263_ VPWR VGND _07274_ sg13g2_a21oi_1
X_27013_ _04635_ _07271_ _07274_ VPWR VGND _07275_ sg13g2_a21oi_1
X_27014_ _12095_ _07267_ _07268_ _07275_ VPWR VGND 
+ _07276_
+ sg13g2_nor4_1
X_27015_ _07256_ _07266_ _07276_ VPWR VGND _07277_ sg13g2_nor3_1
X_27016_ _07277_ _05483_ VPWR VGND _07278_ sg13g2_nand2b_1
X_27017_ _07173_ _07182_ _07246_ _07278_ VPWR VGND 
+ _07279_
+ sg13g2_a22oi_1
X_27018_ \atbs_core_0.spike_memory_0.n2361_o[9]\ _04373_ VPWR VGND _07280_ sg13g2_nor2_1
X_27019_ \atbs_core_0.spike_memory_0.n2358_o[9]\ _04606_ VPWR VGND _07281_ sg13g2_nor2_1
X_27020_ _04513_ _02125_ VPWR VGND _07282_ sg13g2_nor2_1
X_27021_ _02292_ _04716_ VPWR VGND _07283_ sg13g2_nor2_1
X_27022_ _04511_ _07282_ _07283_ _04613_ VPWR VGND 
+ _07284_
+ sg13g2_a22oi_1
X_27023_ _02125_ _04518_ VPWR VGND _07285_ sg13g2_nand2b_1
X_27024_ _03984_ _02292_ _07285_ VPWR VGND _07286_ sg13g2_o21ai_1
X_27025_ _04517_ _07286_ _04521_ VPWR VGND _07287_ sg13g2_a21oi_1
X_27026_ _04608_ _07284_ _07287_ VPWR VGND _07288_ sg13g2_a21oi_1
X_27027_ _04505_ _07280_ _07281_ _07288_ VPWR VGND 
+ _07289_
+ sg13g2_nor4_1
X_27028_ \atbs_core_0.spike_memory_0.n2369_o[9]\ _04525_ VPWR VGND _07290_ sg13g2_nor2_1
X_27029_ \atbs_core_0.spike_memory_0.n2366_o[9]\ _04549_ VPWR VGND _07291_ sg13g2_nor2_1
X_27030_ _04553_ _02035_ VPWR VGND _07292_ sg13g2_nor2_1
X_27031_ _02056_ _04555_ VPWR VGND _07293_ sg13g2_nor2_1
X_27032_ _04531_ _07292_ _07293_ _04557_ VPWR VGND 
+ _07294_
+ sg13g2_a22oi_1
X_27033_ _02035_ _04559_ VPWR VGND _07295_ sg13g2_nand2b_1
X_27034_ _04539_ _02056_ _07295_ VPWR VGND _07296_ sg13g2_o21ai_1
X_27035_ _04538_ _07296_ _04562_ VPWR VGND _07297_ sg13g2_a21oi_1
X_27036_ _04551_ _07294_ _07297_ VPWR VGND _07298_ sg13g2_a21oi_1
X_27037_ _04604_ _07290_ _07291_ _07298_ VPWR VGND 
+ _07299_
+ sg13g2_nor4_1
X_27038_ _03925_ _07289_ _07299_ VPWR VGND _07300_ sg13g2_nor3_1
X_27039_ \atbs_core_0.spike_memory_0.n2365_o[9]\ _04506_ VPWR VGND _07301_ sg13g2_nor2_1
X_27040_ \atbs_core_0.spike_memory_0.n2362_o[9]\ _04508_ VPWR VGND _07302_ sg13g2_nor2_1
X_27041_ _04535_ _12563_ VPWR VGND _07303_ sg13g2_nor2_1
X_27042_ _02009_ _04555_ VPWR VGND _07304_ sg13g2_nor2_1
X_27043_ _04378_ _07303_ _07304_ _04384_ VPWR VGND 
+ _07305_
+ sg13g2_a22oi_1
X_27044_ _12563_ _05544_ VPWR VGND _07306_ sg13g2_nand2b_1
X_27045_ _03755_ _02009_ _07306_ VPWR VGND _07307_ sg13g2_o21ai_1
X_27046_ _04388_ _07307_ _04393_ VPWR VGND _07308_ sg13g2_a21oi_1
X_27047_ _04377_ _07305_ _07308_ VPWR VGND _07309_ sg13g2_a21oi_1
X_27048_ _03968_ _07301_ _07302_ _07309_ VPWR VGND 
+ _07310_
+ sg13g2_nor4_1
X_27049_ \atbs_core_0.spike_memory_0.n2373_o[9]\ _12088_ VPWR VGND _07311_ sg13g2_nor2_1
X_27050_ \atbs_core_0.spike_memory_0.n2370_o[9]\ _04528_ VPWR VGND _07312_ sg13g2_nor2_1
X_27051_ _03934_ _02090_ VPWR VGND _07313_ sg13g2_nor2_1
X_27052_ _02113_ _04570_ VPWR VGND _07314_ sg13g2_nor2_1
X_27053_ _04568_ _07313_ _07314_ _04536_ VPWR VGND 
+ _07315_
+ sg13g2_a22oi_1
X_27054_ _02090_ _04361_ VPWR VGND _07316_ sg13g2_nand2b_1
X_27055_ _04574_ _02113_ _07316_ VPWR VGND _07317_ sg13g2_o21ai_1
X_27056_ _04573_ _07317_ _04542_ VPWR VGND _07318_ sg13g2_a21oi_1
X_27057_ _04530_ _07315_ _07318_ VPWR VGND _07319_ sg13g2_a21oi_1
X_27058_ _04126_ _07311_ _07312_ _07319_ VPWR VGND 
+ _07320_
+ sg13g2_nor4_1
X_27059_ _04547_ _07310_ _07320_ VPWR VGND _07321_ sg13g2_nor3_1
X_27060_ _07549_ _07300_ _07321_ VPWR VGND _07322_ sg13g2_nor3_1
X_27061_ _04503_ _07279_ _07322_ VPWR VGND \atbs_core_0.spike_memory_0.n2550_o[9]\ sg13g2_a21o_1
X_27062_ _08518_ _08891_ _08489_ VPWR VGND _07323_ sg13g2_nand3_1
X_27063_ _08486_ _07323_ VPWR VGND _07324_ sg13g2_nor2_1
X_27064_ _08878_ _08882_ _07324_ VPWR VGND _07325_ sg13g2_nand3_1
X_27065_ _08907_ _07325_ VPWR VGND _07326_ sg13g2_or2_1
X_27066_ _07326_ VPWR VGND _07327_ sg13g2_buf_1
X_27067_ _12416_ _07327_ VPWR VGND _07328_ sg13g2_nor2_1
X_27068_ _10586_ _12404_ _07328_ VPWR VGND _07329_ sg13g2_nand3_1
X_27069_ _08860_ _07329_ VPWR VGND _07330_ sg13g2_nor2_1
X_27070_ _08854_ _12415_ _07330_ VPWR VGND _07331_ sg13g2_nand3_1
X_27071_ _12443_ _07331_ VPWR VGND _07332_ sg13g2_nor2_1
X_27072_ _08943_ _12449_ _07332_ VPWR VGND _07333_ sg13g2_nand3_1
X_27073_ _07333_ VPWR VGND _07334_ sg13g2_buf_1
X_27074_ _08762_ _09035_ _07334_ VPWR VGND \atbs_core_0.time_measurement_0.n2214_o\ sg13g2_nor3_1
X_27075_ \atbs_core_0.time_measurement_0.n2214_o\ _00022_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[0]\ sg13g2_nor2b_1
X_27076_ _09048_ _07329_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[10]\ sg13g2_xnor2_1
X_27077_ _12415_ _07330_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[11]\ sg13g2_xor2_1
X_27078_ _12415_ _07330_ VPWR VGND _07335_ sg13g2_nand2_1
X_27079_ _08854_ _07335_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[12]\ sg13g2_xnor2_1
X_27080_ _12435_ _07331_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[13]\ sg13g2_xnor2_1
X_27081_ _09868_ _07332_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[14]\ sg13g2_xnor2_1
X_27082_ _08943_ _07332_ VPWR VGND _07336_ sg13g2_nand2_1
X_27083_ _12449_ _07336_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[15]\ sg13g2_xnor2_1
X_27084_ _08729_ _07334_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[16]\ sg13g2_xnor2_1
X_27085_ _09035_ _07334_ VPWR VGND _07337_ sg13g2_nor2_1
X_27086_ _08762_ _07337_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[17]\ sg13g2_xnor2_1
X_27087_ _08894_ _08892_ VPWR VGND _07338_ sg13g2_nand2_1
X_27088_ _08888_ _07338_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[2]\ sg13g2_xnor2_1
X_27089_ _08885_ _07323_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[3]\ sg13g2_xnor2_1
X_27090_ _08884_ _07324_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[4]\ sg13g2_xnor2_1
X_27091_ _08883_ _07324_ VPWR VGND _07339_ sg13g2_nand2_1
X_27092_ _08879_ _07339_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[5]\ sg13g2_xnor2_1
X_27093_ _08557_ _07325_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[6]\ sg13g2_xnor2_1
X_27094_ _12400_ _07327_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[7]\ sg13g2_xnor2_1
X_27095_ _10586_ _07328_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[8]\ sg13g2_xor2_1
X_27096_ _10586_ _07328_ VPWR VGND _07340_ sg13g2_nand2_1
X_27097_ _12404_ _07340_ VPWR VGND \atbs_core_0.time_measurement_0.n2218_o[9]\ sg13g2_xnor2_1
X_27098_ _07617_ _07575_ VPWR VGND _07341_ sg13g2_nor2_1
X_27099_ _07578_ VPWR VGND _07342_ sg13g2_inv_1
X_27100_ _07577_ VPWR VGND _07343_ sg13g2_inv_1
X_27101_ _07586_ _07596_ VPWR VGND _07344_ sg13g2_nor2_1
X_27102_ _07585_ _07344_ VPWR VGND _07345_ sg13g2_nor2_1
X_27103_ _07343_ _07578_ _07596_ _07586_ _07345_ VPWR 
+ VGND
+ _07346_ sg13g2_a221oi_1
X_27104_ _07577_ _07342_ _07346_ VPWR VGND _07347_ sg13g2_a21oi_1
X_27105_ _07587_ _07347_ VPWR VGND _07348_ sg13g2_nand2_1
X_27106_ _07587_ _07347_ _07622_ VPWR VGND _07349_ sg13g2_o21ai_1
X_27107_ _07592_ _07348_ _07349_ VPWR VGND _07350_ sg13g2_nand3_1
X_27108_ _07593_ _07350_ VPWR VGND _07351_ sg13g2_and2_1
X_27109_ _07581_ _07351_ _12205_ VPWR VGND _07352_ sg13g2_a21o_1
X_27110_ _07581_ _07351_ _07352_ VPWR VGND _07353_ sg13g2_o21ai_1
X_27111_ _07617_ _07575_ _07571_ VPWR VGND _07354_ sg13g2_a21oi_1
X_27112_ _07341_ _07353_ _07354_ VPWR VGND _07355_ sg13g2_o21ai_1
X_27113_ _12205_ _07582_ _07572_ _07355_ VPWR VGND 
+ _07356_
+ sg13g2_a22oi_1
X_27114_ _12205_ _07582_ VPWR VGND _07357_ sg13g2_nor2_1
X_27115_ _07675_ VPWR VGND _07358_ sg13g2_inv_1
X_27116_ _07356_ _07357_ _07358_ VPWR VGND _07359_ sg13g2_o21ai_1
X_27117_ _07359_ VPWR VGND _07360_ sg13g2_buf_1
X_27118_ _07594_ _07360_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[0]\ sg13g2_nor2_1
X_27119_ _07594_ _07586_ VPWR VGND _07361_ sg13g2_xnor2_1
X_27120_ _07360_ _07361_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[1]\ sg13g2_nor2_1
X_27121_ _07594_ _07586_ VPWR VGND _07362_ sg13g2_nand2_1
X_27122_ _07342_ _07362_ VPWR VGND _07363_ sg13g2_xnor2_1
X_27123_ _07360_ _07363_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[2]\ sg13g2_nor2_1
X_27124_ _07587_ VPWR VGND _07364_ sg13g2_inv_1
X_27125_ _07594_ _07586_ _07578_ VPWR VGND _07365_ sg13g2_nand3_1
X_27126_ _07364_ _07365_ VPWR VGND _07366_ sg13g2_xnor2_1
X_27127_ _07360_ _07366_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[3]\ sg13g2_nor2_1
X_27128_ _07364_ _07365_ VPWR VGND _07367_ sg13g2_nor2_1
X_27129_ _07591_ _07367_ VPWR VGND _07368_ sg13g2_xnor2_1
X_27130_ _07360_ _07368_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[4]\ sg13g2_nor2_1
X_27131_ _07591_ _07367_ VPWR VGND _07369_ sg13g2_nand2_1
X_27132_ _07581_ _07369_ VPWR VGND _07370_ sg13g2_xor2_1
X_27133_ _07360_ _07370_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[5]\ sg13g2_nor2_1
X_27134_ _07591_ _07581_ _07367_ VPWR VGND _07371_ sg13g2_nand3_1
X_27135_ _07575_ _07371_ VPWR VGND _07372_ sg13g2_xor2_1
X_27136_ _07360_ _07372_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[6]\ sg13g2_nor2_1
X_27137_ _07591_ _07581_ _07575_ _07367_ VPWR VGND 
+ _07373_
+ sg13g2_nand4_1
X_27138_ _07570_ _07373_ VPWR VGND _07374_ sg13g2_xnor2_1
X_27139_ _07360_ _07374_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[7]\ sg13g2_nor2_1
X_27140_ _07570_ _07373_ VPWR VGND _07375_ sg13g2_nor2_1
X_27141_ _00057_ _07375_ VPWR VGND _07376_ sg13g2_xnor2_1
X_27142_ _07360_ _07376_ VPWR VGND \atbs_core_0.uart_0.uart_rx_0.n3401_o[8]\ sg13g2_nor2b_1
X_27143_ _07660_ _02959_ VPWR VGND _07377_ sg13g2_nand2_1
X_27144_ _07567_ _07675_ _07608_ _07377_ VPWR VGND 
+ \atbs_core_0.uart_0.uart_rx_0.n3445_o\
+ sg13g2_nor4_1
X_27145_ _07611_ VPWR VGND _07378_ sg13g2_inv_1
X_27146_ _07580_ _07378_ VPWR VGND _07379_ sg13g2_nand2_1
X_27147_ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[7]\ VPWR VGND _07380_ sg13g2_inv_1
X_27148_ _07343_ _07625_ VPWR VGND _07381_ sg13g2_nor2_1
X_27149_ _07622_ _07623_ _07625_ _07343_ VPWR VGND 
+ _07382_
+ sg13g2_a22oi_1
X_27150_ _07381_ _07382_ _07628_ VPWR VGND _07383_ sg13g2_o21ai_1
X_27151_ _07630_ _07383_ _07622_ VPWR VGND _07384_ sg13g2_a21o_1
X_27152_ _07630_ _07383_ _07384_ VPWR VGND _07385_ sg13g2_o21ai_1
X_27153_ _07632_ _07590_ VPWR VGND _07386_ sg13g2_nor2b_1
X_27154_ _07633_ _07385_ _07386_ VPWR VGND _07387_ sg13g2_a21oi_1
X_27155_ _07610_ _07387_ VPWR VGND _07388_ sg13g2_nor2_1
X_27156_ _07610_ _07387_ _12205_ VPWR VGND _07389_ sg13g2_a21oi_1
X_27157_ _07388_ _07389_ VPWR VGND _07390_ sg13g2_nor2_1
X_27158_ _07620_ _07390_ VPWR VGND _07391_ sg13g2_nand2_1
X_27159_ _07619_ _07391_ VPWR VGND _07392_ sg13g2_and2_1
X_27160_ _07380_ _07392_ VPWR VGND _07393_ sg13g2_nand2_1
X_27161_ _07380_ _07392_ _07569_ VPWR VGND _07394_ sg13g2_o21ai_1
X_27162_ _07379_ _07393_ _07394_ VPWR VGND _07395_ sg13g2_nand3_1
X_27163_ _07580_ _07378_ _07395_ VPWR VGND _07396_ sg13g2_o21ai_1
X_27164_ _07396_ VPWR VGND _07397_ sg13g2_buf_1
X_27165_ _07615_ _07397_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[0]\ sg13g2_nor2_1
X_27166_ _07615_ _07623_ VPWR VGND _07398_ sg13g2_xnor2_1
X_27167_ _07397_ _07398_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[1]\ sg13g2_nor2_1
X_27168_ _07615_ _07623_ VPWR VGND _07399_ sg13g2_nand2_1
X_27169_ _07625_ _07399_ VPWR VGND _07400_ sg13g2_xor2_1
X_27170_ _07397_ _07400_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[2]\ sg13g2_nor2_1
X_27171_ _07630_ VPWR VGND _07401_ sg13g2_inv_1
X_27172_ _07615_ _07623_ _07625_ VPWR VGND _07402_ sg13g2_nand3_1
X_27173_ _07401_ _07402_ VPWR VGND _07403_ sg13g2_xnor2_1
X_27174_ _07397_ _07403_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[3]\ sg13g2_nor2_1
X_27175_ _07401_ _07402_ VPWR VGND _07404_ sg13g2_nor2_1
X_27176_ _07632_ _07404_ VPWR VGND _07405_ sg13g2_xnor2_1
X_27177_ _07397_ _07405_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[4]\ sg13g2_nor2_1
X_27178_ _07632_ _07404_ VPWR VGND _07406_ sg13g2_nand2_1
X_27179_ _07610_ _07406_ VPWR VGND _07407_ sg13g2_xor2_1
X_27180_ _07397_ _07407_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[5]\ sg13g2_nor2_1
X_27181_ _07610_ _07632_ _07404_ VPWR VGND _07408_ sg13g2_nand3_1
X_27182_ _07618_ _07408_ VPWR VGND _07409_ sg13g2_xor2_1
X_27183_ _07397_ _07409_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[6]\ sg13g2_nor2_1
X_27184_ _07618_ _07610_ _07632_ _07404_ VPWR VGND 
+ _07410_
+ sg13g2_nand4_1
X_27185_ _07380_ _07410_ VPWR VGND _07411_ sg13g2_xnor2_1
X_27186_ _07397_ _07411_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[7]\ sg13g2_nor2_1
X_27187_ _07380_ _07410_ VPWR VGND _07412_ sg13g2_nor2_1
X_27188_ _07611_ _07412_ VPWR VGND _07413_ sg13g2_xnor2_1
X_27189_ _07397_ _07413_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3277_o[8]\ sg13g2_nor2_1
X_27190_ _07647_ _07642_ VPWR VGND _07414_ sg13g2_nor2_1
X_27191_ _02961_ _07414_ VPWR VGND \atbs_core_0.uart_0.uart_tx_0.n3341_o\ sg13g2_and2_1
X_27192_ _12308_ VPWR VGND _07415_ sg13g2_inv_1
X_27193_ _07415_ _12303_ _12300_ VPWR VGND _07416_ sg13g2_a21oi_1
X_27194_ _07415_ _12303_ VPWR VGND _07417_ sg13g2_nor2_1
X_27195_ _12307_ _12163_ VPWR VGND _07418_ sg13g2_nand2_1
X_27196_ _07416_ _07417_ _07418_ VPWR VGND _07419_ sg13g2_o21ai_1
X_27197_ _12307_ _12162_ VPWR VGND _07420_ sg13g2_nand2b_1
X_27198_ _07419_ _07420_ _12316_ VPWR VGND phi_bias_1_o sg13g2_a21oi_1
X_27199_ _12307_ _12305_ _12316_ VPWR VGND _07421_ sg13g2_o21ai_1
X_27200_ _12162_ _12305_ VPWR VGND _07422_ sg13g2_xor2_1
X_27201_ _12300_ _07422_ VPWR VGND _07423_ sg13g2_nand2_1
X_27202_ _12315_ _07418_ _07423_ VPWR VGND _07424_ sg13g2_nand3_1
X_27203_ _12162_ _12305_ _12308_ VPWR VGND _07425_ sg13g2_o21ai_1
X_27204_ _12308_ _07424_ _07425_ VPWR VGND _07426_ sg13g2_o21ai_1
X_27205_ _12162_ _12315_ VPWR VGND _07427_ sg13g2_xor2_1
X_27206_ _12308_ _12305_ VPWR VGND _07428_ sg13g2_xor2_1
X_27207_ _12300_ _12301_ _07427_ _07428_ VPWR VGND 
+ _07429_
+ sg13g2_nand4_1
X_27208_ _12308_ _12305_ VPWR VGND _07430_ sg13g2_nor2_1
X_27209_ _12163_ \atbs_core_0.sc_noc_generator_1.counter_value[7]\ _07427_ _07430_ VPWR VGND 
+ _07431_
+ sg13g2_a22oi_1
X_27210_ _12300_ _07415_ _12162_ _12305_ VPWR VGND 
+ _07432_
+ sg13g2_nor4_1
X_27211_ _12308_ _07423_ VPWR VGND _07433_ sg13g2_nor2_1
X_27212_ _07432_ _07433_ _12315_ VPWR VGND _07434_ sg13g2_o21ai_1
X_27213_ _12300_ VPWR VGND _07435_ sg13g2_inv_1
X_27214_ _07435_ _12308_ _12162_ _12305_ VPWR VGND 
+ _07436_
+ sg13g2_nand4_1
X_27215_ _07434_ _07436_ VPWR VGND _07437_ sg13g2_nand2_1
X_27216_ _12293_ \atbs_core_0.sc_noc_generator_1.counter_value[3]\ _12295_ \atbs_core_0.sc_noc_generator_1.counter_value[4]\ VPWR VGND 
+ _07438_
+ sg13g2_nor4_1
X_27217_ _07437_ _07438_ VPWR VGND _07439_ sg13g2_nand2_1
X_27218_ _07439_ _07429_ _12292_ VPWR VGND _07440_ sg13g2_a21oi_1
X_27219_ _07429_ _07431_ _07440_ VPWR VGND _07441_ sg13g2_a21oi_1
X_27220_ _07421_ _07426_ _07441_ VPWR VGND phi_bias_2_o sg13g2_a21oi_1
X_27221_ _12333_ _12338_ VPWR VGND _07442_ sg13g2_nand2_1
X_27222_ _12340_ VPWR VGND _07443_ sg13g2_inv_1
X_27223_ _07443_ _12331_ _12329_ VPWR VGND _07444_ sg13g2_a21o_1
X_27224_ _07443_ _12331_ _07444_ VPWR VGND _07445_ sg13g2_o21ai_1
X_27225_ _12333_ _12338_ VPWR VGND _07446_ sg13g2_nor2_1
X_27226_ _07442_ _07445_ _07446_ VPWR VGND _07447_ sg13g2_a21oi_1
X_27227_ _12346_ _07447_ VPWR VGND phi_cmfb_1_o sg13g2_nor2_1
X_27228_ _12169_ _12334_ VPWR VGND _07448_ sg13g2_nor2_1
X_27229_ _12169_ _12334_ VPWR VGND _07449_ sg13g2_xor2_1
X_27230_ _12340_ _12329_ VPWR VGND _07450_ sg13g2_nor2b_1
X_27231_ _12340_ _07448_ _07449_ _07450_ VPWR VGND 
+ _07451_
+ sg13g2_a22oi_1
X_27232_ _12340_ _12169_ _12334_ VPWR VGND _07452_ sg13g2_nand3_1
X_27233_ _07451_ _07452_ _12346_ VPWR VGND _07453_ sg13g2_mux2_1
X_27234_ _12322_ _12321_ \atbs_core_0.sc_noc_generator_2.counter_value[3]\ _12324_ VPWR VGND 
+ _07454_
+ sg13g2_nor4_1
X_27235_ _12329_ _12340_ \atbs_core_0.sc_noc_generator_2.counter_value[4]\ VPWR VGND _07455_ sg13g2_a21oi_1
X_27236_ _07454_ _07455_ VPWR VGND _07456_ sg13g2_nand2_1
X_27237_ _12334_ _12347_ _12340_ VPWR VGND _07457_ sg13g2_o21ai_1
X_27238_ _12334_ _12347_ VPWR VGND _07458_ sg13g2_nand2_1
X_27239_ _07457_ _07458_ _12337_ VPWR VGND _07459_ sg13g2_a21oi_1
X_27240_ _12340_ _12169_ _12345_ VPWR VGND _07460_ sg13g2_a21oi_1
X_27241_ _12340_ _12169_ _12345_ VPWR VGND _07461_ sg13g2_o21ai_1
X_27242_ _12333_ _07460_ _07461_ VPWR VGND _07462_ sg13g2_o21ai_1
X_27243_ _07453_ _07462_ VPWR VGND _07463_ sg13g2_nand2_1
X_27244_ _12339_ _07459_ _07463_ VPWR VGND _07464_ sg13g2_o21ai_1
X_27245_ _07453_ _07456_ _07464_ VPWR VGND phi_cmfb_2_o sg13g2_o21ai_1
X_27246_ \atbs_core_0.analog_trigger_0.counter_value[2]\ _11355_ _11353_ \atbs_core_0.analog_trigger_0.counter_value[6]\ VPWR VGND 
+ _07465_
+ sg13g2_or4_1
X_27247_ \atbs_core_0.analog_trigger_0.counter_value[1]\ _11345_ _11351_ _07465_ VPWR VGND 
+ phi_comp_o
+ sg13g2_nor4_1
X_27248_ \atbs_core_0.dac_control_1.n2062_o\ \atbs_core_0.clear_dac\ _07844_ VPWR VGND phi_dac_lower_o sg13g2_and3_1
X_27249_ \atbs_core_0.dac_control_0.n1913_o\ \atbs_core_0.clear_dac\ _07844_ VPWR VGND phi_dac_upper_o sg13g2_and3_1
X_27250_ _12352_ _12354_ _12359_ VPWR VGND _07466_ sg13g2_nand3_1
X_27251_ _12182_ _12362_ _07466_ VPWR VGND _07467_ sg13g2_nor3_1
X_27252_ _12362_ _07466_ _12182_ VPWR VGND _07468_ sg13g2_o21ai_1
X_27253_ _12353_ _07467_ _07468_ VPWR VGND _07469_ sg13g2_o21ai_1
X_27254_ _00029_ _07469_ VPWR VGND phi_res_1_o sg13g2_and2_1
X_27255_ _12354_ _12359_ VPWR VGND _07470_ sg13g2_nand2_1
X_27256_ _00028_ _07470_ VPWR VGND _07471_ sg13g2_nor2_1
X_27257_ _12182_ _12362_ VPWR VGND _07472_ sg13g2_nand2_1
X_27258_ _12182_ _12362_ _07471_ VPWR VGND _07473_ sg13g2_nor3_1
X_27259_ _12352_ _12381_ VPWR VGND _07474_ sg13g2_nor2_1
X_27260_ _07473_ _07474_ _12353_ VPWR VGND _07475_ sg13g2_o21ai_1
X_27261_ _07471_ _07472_ _07475_ VPWR VGND phi_res_2_o sg13g2_o21ai_1
X_27262_ _12279_ VPWR VGND _07476_ sg13g2_inv_1
X_27263_ _07476_ _12274_ _12271_ VPWR VGND _07477_ sg13g2_a21oi_1
X_27264_ _07476_ _12274_ VPWR VGND _07478_ sg13g2_nor2_1
X_27265_ _12278_ _12151_ VPWR VGND _07479_ sg13g2_nand2_1
X_27266_ _07477_ _07478_ _07479_ VPWR VGND _07480_ sg13g2_o21ai_1
X_27267_ _12278_ _12150_ VPWR VGND _07481_ sg13g2_nand2b_1
X_27268_ _07480_ _07481_ _12287_ VPWR VGND phi_vcm_generator_1_o sg13g2_a21oi_1
X_27269_ _12278_ _12276_ _12287_ VPWR VGND _07482_ sg13g2_o21ai_1
X_27270_ _12150_ _12276_ VPWR VGND _07483_ sg13g2_xor2_1
X_27271_ _12271_ _07483_ VPWR VGND _07484_ sg13g2_nand2_1
X_27272_ _12286_ _07479_ _07484_ VPWR VGND _07485_ sg13g2_nand3_1
X_27273_ _12150_ _12276_ _12279_ VPWR VGND _07486_ sg13g2_o21ai_1
X_27274_ _12279_ _07485_ _07486_ VPWR VGND _07487_ sg13g2_o21ai_1
X_27275_ _12264_ _12263_ _12266_ \atbs_core_0.sc_noc_generator_0.counter_value[3]\ VPWR VGND 
+ _07488_
+ sg13g2_nor4_1
X_27276_ _12271_ _12279_ VPWR VGND _07489_ sg13g2_nand2b_1
X_27277_ _12150_ _12276_ VPWR VGND _07490_ sg13g2_nand2_1
X_27278_ _12150_ _12276_ _07489_ VPWR VGND _07491_ sg13g2_nor3_1
X_27279_ _12279_ _07484_ VPWR VGND _07492_ sg13g2_nor2_1
X_27280_ _07491_ _07492_ _12286_ VPWR VGND _07493_ sg13g2_o21ai_1
X_27281_ _07489_ _07490_ _07493_ VPWR VGND _07494_ sg13g2_o21ai_1
X_27282_ \atbs_core_0.sc_noc_generator_0.counter_value[4]\ _07488_ _07494_ VPWR VGND _07495_ sg13g2_nand3b_1
X_27283_ _12279_ _12276_ VPWR VGND _07496_ sg13g2_xor2_1
X_27284_ _12150_ _12286_ VPWR VGND _07497_ sg13g2_xor2_1
X_27285_ _12271_ _12272_ _07496_ _07497_ VPWR VGND 
+ _07498_
+ sg13g2_nand4_1
X_27286_ _12279_ _12276_ VPWR VGND _07499_ sg13g2_nor2_1
X_27287_ _12151_ \atbs_core_0.sc_noc_generator_0.counter_value[7]\ _07497_ _07499_ VPWR VGND 
+ _07500_
+ sg13g2_a22oi_1
X_27288_ _12263_ _07498_ VPWR VGND _07501_ sg13g2_nor2_1
X_27289_ _07498_ _07500_ _07501_ VPWR VGND _07502_ sg13g2_a21oi_1
X_27290_ _07482_ _07487_ _07495_ _07502_ VPWR VGND 
+ phi_vcm_generator_2_o
+ sg13g2_a22oi_1
X_27291_ \atbs_core_0.n1402_q[0]\ bio_amp_en_o VPWR VGND select_cap_o[0] sg13g2_and2_1
X_27292_ \atbs_core_0.n1402_q[1]\ bio_amp_en_o VPWR VGND select_cap_o[1] sg13g2_and2_1
X_27293_ \atbs_core_0.n1402_q[2]\ bio_amp_en_o VPWR VGND select_cap_o[2] sg13g2_and2_1
X_27294_ \atbs_core_0.n1418_q\ VPWR VGND _07503_ sg13g2_inv_1
X_27295_ _00039_ _07503_ _07653_ VPWR VGND select_spdt_o sg13g2_mux2_1
X_27296_ _07638_ _07649_ VPWR VGND _07504_ sg13g2_xnor2_1
X_27297_ _07638_ _00061_ VPWR VGND _07505_ sg13g2_nor2b_1
X_27298_ _07636_ _07505_ _07640_ VPWR VGND _07506_ sg13g2_nand3b_1
X_27299_ _07640_ _07504_ _07506_ VPWR VGND _07507_ sg13g2_o21ai_1
X_27300_ \atbs_core_0.uart_0.uart_tx_0.n3349_o\ \atbs_core_0.uart_0.uart_tx_0.n3353_o\ \atbs_core_0.uart_0.uart_tx_0.n3351_o\ \atbs_core_0.uart_0.uart_tx_0.n3355_o\ _07645_ _07643_ 
+ VPWR
+ VGND _07508_ sg13g2_mux4_1
X_27301_ \atbs_core_0.uart_0.uart_tx_0.n3348_o\ \atbs_core_0.uart_0.uart_tx_0.n3352_o\ \atbs_core_0.uart_0.uart_tx_0.n3350_o\ \atbs_core_0.uart_0.uart_tx_0.n3354_o\ _07645_ _07643_ 
+ VPWR
+ VGND _07509_ sg13g2_mux4_1
X_27302_ _07644_ _07509_ VPWR VGND _07510_ sg13g2_nor2b_1
X_27303_ _07644_ _07508_ _07510_ VPWR VGND _07511_ sg13g2_a21oi_1
X_27304_ _07640_ _07511_ VPWR VGND _07512_ sg13g2_nor2_1
X_27305_ _07845_ _07507_ _07512_ VPWR VGND _07513_ sg13g2_a21oi_1
X_27306_ _07640_ _07642_ _07647_ VPWR VGND _07514_ sg13g2_a21oi_1
X_27307_ _07505_ _07514_ _07511_ VPWR VGND _07515_ sg13g2_a21o_1
X_27308_ _07642_ _07513_ _07515_ VPWR VGND uart_tx_o sg13g2_o21ai_1
X_27309_ _14577_ VPWR VGND sg13g2_tiehi
X\atbs_core_0.adaptive_ctrl_0.n1778_q$_DFFE_PP0P_  clock_i _00191_ \atbs_core_0.adaptive_ctrl_0.adapt_on_overflow\ _00051_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1779_q$_DFFE_PP0P_  clock_i _00192_ \atbs_core_0.adaptive_ctrl_0.is_empty_interval\ _14571_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1780_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1682_o\ \atbs_core_0.adaptive_ctrl_0.adaptive_strb\ _00054_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1781_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1685_o\ \atbs_core_0.adaptive_ctrl_0.n1781_q\ _00052_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1782_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1689_o\ \atbs_core_0.adaptive_ctrl_0.delta_steps_strb\ _14570_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[0]$_DFFE_PP1P_  clock_i _00193_ _00151_ \atbs_core_0.adaptive_ctrl_0.delta_steps[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[1]$_DFFE_PP0P_  clock_i _00194_ \atbs_core_0.adaptive_ctrl_0.delta_steps[1]\ _00080_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[2]$_DFFE_PP0P_  clock_i _00195_ \atbs_core_0.adaptive_ctrl_0.delta_steps[2]\ _00084_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[3]$_DFFE_PP0P_  clock_i _00196_ \atbs_core_0.adaptive_ctrl_0.delta_steps[3]\ _00082_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[4]$_DFFE_PP0P_  clock_i _00197_ \atbs_core_0.adaptive_ctrl_0.delta_steps[4]\ _00088_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[5]$_DFFE_PP0P_  clock_i _00198_ \atbs_core_0.adaptive_ctrl_0.delta_steps[5]\ _00086_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1783_q[6]$_DFFE_PP0P_  clock_i _00199_ \atbs_core_0.adaptive_ctrl_0.delta_steps[6]\ _00090_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[0]$_DFFE_PP1P_  clock_i _00200_ _00152_ \atbs_core_0.adaptive_ctrl_0.n1784_q[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[1]$_DFFE_PP0P_  clock_i _00201_ \atbs_core_0.adaptive_ctrl_0.n1784_q[1]\ _14569_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[2]$_DFFE_PP0P_  clock_i _00202_ \atbs_core_0.adaptive_ctrl_0.n1784_q[2]\ _14568_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[3]$_DFFE_PP0P_  clock_i _00203_ \atbs_core_0.adaptive_ctrl_0.n1784_q[3]\ _14567_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[4]$_DFFE_PP0P_  clock_i _00204_ \atbs_core_0.adaptive_ctrl_0.n1784_q[4]\ _14566_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[5]$_DFFE_PP0P_  clock_i _00205_ \atbs_core_0.adaptive_ctrl_0.n1784_q[5]\ _14565_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1784_q[6]$_DFFE_PP0P_  clock_i _00206_ \atbs_core_0.adaptive_ctrl_0.n1784_q[6]\ _14564_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[0]$_DFFE_PP1P_  clock_i _00207_ _00153_ \atbs_core_0.adaptive_ctrl_0.n1705_o[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[1]$_DFFE_PP0P_  clock_i _00208_ \atbs_core_0.adaptive_ctrl_0.n1705_o[1]\ _00081_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[2]$_DFFE_PP1P_  clock_i _00209_ _00154_ \atbs_core_0.adaptive_ctrl_0.n1705_o[2]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[3]$_DFFE_PP1P_  clock_i _00210_ _00155_ \atbs_core_0.adaptive_ctrl_0.n1705_o[3]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[4]$_DFFE_PP1P_  clock_i _00211_ _00156_ \atbs_core_0.adaptive_ctrl_0.n1705_o[4]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[5]$_DFFE_PP1P_  clock_i _00212_ _00157_ \atbs_core_0.adaptive_ctrl_0.n1705_o[5]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[6]$_DFFE_PP0P_  clock_i _00213_ \atbs_core_0.adaptive_ctrl_0.n1705_o[6]\ _00091_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1785_q[7]$_DFFE_PP0P_  clock_i _00214_ \atbs_core_0.adaptive_ctrl_0.n1785_q[7]\ _00055_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[0]$_DFFE_PP1P_  clock_i _00215_ _00158_ \atbs_core_0.adaptive_ctrl_0.n1710_o[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[1]$_DFFE_PP1P_  clock_i _00216_ _00159_ \atbs_core_0.adaptive_ctrl_0.n1710_o[1]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[2]$_DFFE_PP1P_  clock_i _00217_ _00160_ \atbs_core_0.adaptive_ctrl_0.n1710_o[2]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[3]$_DFFE_PP1P_  clock_i _00218_ _00161_ \atbs_core_0.adaptive_ctrl_0.n1710_o[3]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[4]$_DFFE_PP1P_  clock_i _00219_ _00162_ \atbs_core_0.adaptive_ctrl_0.n1710_o[4]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[5]$_DFFE_PP1P_  clock_i _00220_ _00163_ \atbs_core_0.adaptive_ctrl_0.n1710_o[5]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[6]$_DFFE_PP0P_  clock_i _00221_ \atbs_core_0.adaptive_ctrl_0.n1710_o[6]\ _00092_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.n1786_q[7]$_DFFE_PP0P_  clock_i _00222_ \atbs_core_0.adaptive_ctrl_0.n1786_q[7]\ _14563_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[0]$_DFFE_PP0N_  clock_i _00223_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[0]\ _14562_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[100]$_DFFE_PP0N_  clock_i _00224_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[10]\ _14561_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[101]$_DFFE_PP0N_  clock_i _00225_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[11]\ _14560_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[102]$_DFFE_PP0N_  clock_i _00226_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[12]\ _14559_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[103]$_DFFE_PP0N_  clock_i _00227_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[13]\ _14558_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[104]$_DFFE_PP0N_  clock_i _00228_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[14]\ _14557_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[105]$_DFFE_PP0N_  clock_i _00229_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[15]\ _14556_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[106]$_DFFE_PP0N_  clock_i _00230_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[16]\ _14555_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[107]$_DFFE_PP0N_  clock_i _00231_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[17]\ _14554_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[108]$_DFFE_PP0N_  clock_i _00232_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[114]\ _14553_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[109]$_DFFE_PP0N_  clock_i _00233_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[115]\ _14552_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[10]$_DFFE_PP0N_  clock_i _00234_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[10]\ _14551_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[110]$_DFFE_PP0N_  clock_i _00235_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[116]\ _14550_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[111]$_DFFE_PP0N_  clock_i _00236_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[117]\ _14549_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[112]$_DFFE_PP0N_  clock_i _00237_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[118]\ _14548_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[113]$_DFFE_PP0N_  clock_i _00238_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[119]\ _14547_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[114]$_DFFE_PP0N_  clock_i _00239_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[6]\ _14546_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[115]$_DFFE_PP0N_  clock_i _00240_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[7]\ _14545_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[116]$_DFFE_PP0N_  clock_i _00241_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[8]\ _14544_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[117]$_DFFE_PP0N_  clock_i _00242_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[9]\ _14543_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[118]$_DFFE_PP0N_  clock_i _00243_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[10]\ _14542_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[119]$_DFFE_PP0N_  clock_i _00244_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[11]\ _14541_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[11]$_DFFE_PP0N_  clock_i _00245_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[11]\ _14540_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[120]$_DFFE_PP0N_  clock_i _00246_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[12]\ _14539_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[121]$_DFFE_PP0N_  clock_i _00247_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[13]\ _14538_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[122]$_DFFE_PP0N_  clock_i _00248_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[14]\ _14537_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[123]$_DFFE_PP0N_  clock_i _00249_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[15]\ _14536_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[124]$_DFFE_PP0N_  clock_i _00250_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[16]\ _14535_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[125]$_DFFE_PP0N_  clock_i _00251_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2654_o[17]\ _14534_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[126]$_DFFE_PP0N_  clock_i _00252_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[133]\ _14533_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[127]$_DFFE_PP0N_  clock_i _00253_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[134]\ _14532_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[128]$_DFFE_PP0N_  clock_i _00254_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[135]\ _14531_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[129]$_DFFE_PP0N_  clock_i _00255_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[136]\ _14530_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[12]$_DFFE_PP0N_  clock_i _00256_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[12]\ _14529_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[130]$_DFFE_PP0N_  clock_i _00257_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[137]\ _14528_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[131]$_DFFE_PP0N_  clock_i _00258_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[138]\ _14527_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[132]$_DFFE_PP0N_  clock_i _00259_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[6]\ _14526_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[133]$_DFFE_PP0N_  clock_i _00260_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[7]\ _14525_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[134]$_DFFE_PP0N_  clock_i _00261_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[8]\ _14524_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[135]$_DFFE_PP0N_  clock_i _00262_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[9]\ _14523_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[136]$_DFFE_PP0N_  clock_i _00263_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[10]\ _14522_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[137]$_DFFE_PP0N_  clock_i _00264_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[11]\ _14521_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[138]$_DFFE_PP0N_  clock_i _00265_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[12]\ _14520_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[139]$_DFFE_PP0N_  clock_i _00266_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[13]\ _14519_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[13]$_DFFE_PP0N_  clock_i _00267_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[13]\ _14518_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[140]$_DFFE_PP0N_  clock_i _00268_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[14]\ _14517_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[141]$_DFFE_PP0N_  clock_i _00269_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[15]\ _14516_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[142]$_DFFE_PP0N_  clock_i _00270_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[16]\ _14515_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[143]$_DFFE_PP0N_  clock_i _00271_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2657_o[17]\ _14514_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[144]$_DFFE_PP0N_  clock_i _00272_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[152]\ _14513_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[145]$_DFFE_PP0N_  clock_i _00273_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[153]\ _14512_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[146]$_DFFE_PP0N_  clock_i _00274_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[154]\ _14511_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[147]$_DFFE_PP0N_  clock_i _00275_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[155]\ _14510_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[148]$_DFFE_PP0N_  clock_i _00276_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[156]\ _14509_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[149]$_DFFE_PP0N_  clock_i _00277_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[157]\ _14508_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[14]$_DFFE_PP0N_  clock_i _00278_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[14]\ _14507_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[150]$_DFFE_PP0N_  clock_i _00279_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[6]\ _14506_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[151]$_DFFE_PP0N_  clock_i _00280_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[7]\ _14505_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[152]$_DFFE_PP0N_  clock_i _00281_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[8]\ _14504_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[153]$_DFFE_PP0N_  clock_i _00282_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[9]\ _14503_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[154]$_DFFE_PP0N_  clock_i _00283_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[10]\ _14502_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[155]$_DFFE_PP0N_  clock_i _00284_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[11]\ _14501_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[156]$_DFFE_PP0N_  clock_i _00285_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[12]\ _14500_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[157]$_DFFE_PP0N_  clock_i _00286_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[13]\ _14499_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[158]$_DFFE_PP0N_  clock_i _00287_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[14]\ _14498_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[159]$_DFFE_PP0N_  clock_i _00288_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[15]\ _14497_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[15]$_DFFE_PP0N_  clock_i _00289_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[15]\ _14496_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[160]$_DFFE_PP0N_  clock_i _00290_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[16]\ _14495_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[161]$_DFFE_PP0N_  clock_i _00291_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2660_o[17]\ _14494_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[162]$_DFFE_PP0N_  clock_i _00292_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[171]\ _14493_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[163]$_DFFE_PP0N_  clock_i _00293_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[172]\ _14492_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[164]$_DFFE_PP0N_  clock_i _00294_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[173]\ _14491_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[165]$_DFFE_PP0N_  clock_i _00295_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[174]\ _14490_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[166]$_DFFE_PP0N_  clock_i _00296_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[175]\ _14489_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[167]$_DFFE_PP0N_  clock_i _00297_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[176]\ _14488_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[168]$_DFFE_PP0N_  clock_i _00298_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[6]\ _14487_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[169]$_DFFE_PP0N_  clock_i _00299_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[7]\ _14486_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[16]$_DFFE_PP0N_  clock_i _00300_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[16]\ _14485_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[170]$_DFFE_PP0N_  clock_i _00301_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[8]\ _14484_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[171]$_DFFE_PP0N_  clock_i _00302_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[9]\ _14483_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[172]$_DFFE_PP0N_  clock_i _00303_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[10]\ _14482_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[173]$_DFFE_PP0N_  clock_i _00304_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[11]\ _14481_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[174]$_DFFE_PP0N_  clock_i _00305_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[12]\ _14480_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[175]$_DFFE_PP0N_  clock_i _00306_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[13]\ _14479_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[176]$_DFFE_PP0N_  clock_i _00307_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[14]\ _14478_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[177]$_DFFE_PP0N_  clock_i _00308_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[15]\ _14477_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[178]$_DFFE_PP0N_  clock_i _00309_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[16]\ _14476_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[179]$_DFFE_PP0N_  clock_i _00310_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2663_o[17]\ _14475_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[17]$_DFFE_PP0N_  clock_i _00311_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[17]\ _14474_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[180]$_DFFE_PP0N_  clock_i _00312_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[190]\ _14473_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[181]$_DFFE_PP0N_  clock_i _00313_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[191]\ _14472_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[182]$_DFFE_PP0N_  clock_i _00314_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[192]\ _14471_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[183]$_DFFE_PP0N_  clock_i _00315_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[193]\ _14470_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[184]$_DFFE_PP0N_  clock_i _00316_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[194]\ _14469_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[185]$_DFFE_PP0N_  clock_i _00317_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[195]\ _14468_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[186]$_DFFE_PP0N_  clock_i _00318_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[6]\ _14467_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[187]$_DFFE_PP0N_  clock_i _00319_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[7]\ _14466_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[188]$_DFFE_PP0N_  clock_i _00320_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[8]\ _14465_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[189]$_DFFE_PP0N_  clock_i _00321_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[9]\ _14464_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[18]$_DFFE_PP0N_  clock_i _00322_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[19]\ _14463_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[190]$_DFFE_PP0N_  clock_i _00323_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[10]\ _14462_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[191]$_DFFE_PP0N_  clock_i _00324_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[11]\ _14461_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[192]$_DFFE_PP0N_  clock_i _00325_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[12]\ _14460_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[193]$_DFFE_PP0N_  clock_i _00326_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[13]\ _14459_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[194]$_DFFE_PP0N_  clock_i _00327_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[14]\ _14458_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[195]$_DFFE_PP0N_  clock_i _00328_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[15]\ _14457_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[196]$_DFFE_PP0N_  clock_i _00329_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[16]\ _14456_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[197]$_DFFE_PP0N_  clock_i _00330_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2666_o[17]\ _14455_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[198]$_DFFE_PP0N_  clock_i _00331_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[209]\ _14454_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[199]$_DFFE_PP0N_  clock_i _00332_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[210]\ _14453_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[19]$_DFFE_PP0N_  clock_i _00333_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[20]\ _14452_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[1]$_DFFE_PP0N_  clock_i _00334_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[1]\ _14451_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[200]$_DFFE_PP0N_  clock_i _00335_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[211]\ _14450_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[201]$_DFFE_PP0N_  clock_i _00336_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[212]\ _14449_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[202]$_DFFE_PP0N_  clock_i _00337_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[213]\ _14448_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[203]$_DFFE_PP0N_  clock_i _00338_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[214]\ _14447_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[204]$_DFFE_PP0N_  clock_i _00339_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[6]\ _14446_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[205]$_DFFE_PP0N_  clock_i _00340_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[7]\ _14445_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[206]$_DFFE_PP0N_  clock_i _00341_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[8]\ _14444_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[207]$_DFFE_PP0N_  clock_i _00342_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[9]\ _14443_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[208]$_DFFE_PP0N_  clock_i _00343_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[10]\ _14442_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[209]$_DFFE_PP0N_  clock_i _00344_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[11]\ _14441_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[20]$_DFFE_PP0N_  clock_i _00345_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[21]\ _14440_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[210]$_DFFE_PP0N_  clock_i _00346_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[12]\ _14439_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[211]$_DFFE_PP0N_  clock_i _00347_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[13]\ _14438_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[212]$_DFFE_PP0N_  clock_i _00348_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[14]\ _14437_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[213]$_DFFE_PP0N_  clock_i _00349_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[15]\ _14436_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[214]$_DFFE_PP0N_  clock_i _00350_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[16]\ _14435_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[215]$_DFFE_PP0N_  clock_i _00351_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2669_o[17]\ _14434_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[216]$_DFFE_PP0N_  clock_i _00352_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[228]\ _14433_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[217]$_DFFE_PP0N_  clock_i _00353_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[229]\ _14432_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[218]$_DFFE_PP0N_  clock_i _00354_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[230]\ _14431_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[219]$_DFFE_PP0N_  clock_i _00355_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[231]\ _14430_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[21]$_DFFE_PP0N_  clock_i _00356_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[22]\ _14429_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[220]$_DFFE_PP0N_  clock_i _00357_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[232]\ _14428_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[221]$_DFFE_PP0N_  clock_i _00358_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[233]\ _14427_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[222]$_DFFE_PP0N_  clock_i _00359_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[6]\ _14426_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[223]$_DFFE_PP0N_  clock_i _00360_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[7]\ _14425_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[224]$_DFFE_PP0N_  clock_i _00361_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[8]\ _14424_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[225]$_DFFE_PP0N_  clock_i _00362_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[9]\ _14423_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[226]$_DFFE_PP0N_  clock_i _00363_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[10]\ _14422_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[227]$_DFFE_PP0N_  clock_i _00364_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[11]\ _14421_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[228]$_DFFE_PP0N_  clock_i _00365_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[12]\ _14420_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[229]$_DFFE_PP0N_  clock_i _00366_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[13]\ _14419_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[22]$_DFFE_PP0N_  clock_i _00367_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[23]\ _14418_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[230]$_DFFE_PP0N_  clock_i _00368_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[14]\ _14417_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[231]$_DFFE_PP0N_  clock_i _00369_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[15]\ _14416_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[232]$_DFFE_PP0N_  clock_i _00370_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[16]\ _14415_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[233]$_DFFE_PP0N_  clock_i _00371_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2672_o[17]\ _14414_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[234]$_DFFE_PP0N_  clock_i _00372_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[247]\ _14413_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[235]$_DFFE_PP0N_  clock_i _00373_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[248]\ _14412_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[236]$_DFFE_PP0N_  clock_i _00374_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[249]\ _14411_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[237]$_DFFE_PP0N_  clock_i _00375_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[250]\ _14410_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[238]$_DFFE_PP0N_  clock_i _00376_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[251]\ _14409_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[239]$_DFFE_PP0N_  clock_i _00377_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[252]\ _14408_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[23]$_DFFE_PP0N_  clock_i _00378_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[24]\ _14407_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[240]$_DFFE_PP0N_  clock_i _00379_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[6]\ _14406_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[241]$_DFFE_PP0N_  clock_i _00380_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[7]\ _14405_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[242]$_DFFE_PP0N_  clock_i _00381_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[8]\ _14404_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[243]$_DFFE_PP0N_  clock_i _00382_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[9]\ _14403_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[244]$_DFFE_PP0N_  clock_i _00383_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[10]\ _14402_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[245]$_DFFE_PP0N_  clock_i _00384_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[11]\ _14401_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[246]$_DFFE_PP0N_  clock_i _00385_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[12]\ _14400_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[247]$_DFFE_PP0N_  clock_i _00386_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[13]\ _14399_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[248]$_DFFE_PP0N_  clock_i _00387_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[14]\ _14398_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[249]$_DFFE_PP0N_  clock_i _00388_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[15]\ _14397_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[24]$_DFFE_PP0N_  clock_i _00389_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[6]\ _14396_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[250]$_DFFE_PP0N_  clock_i _00390_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[16]\ _14395_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[251]$_DFFE_PP0N_  clock_i _00391_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2675_o[17]\ _14394_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[252]$_DFFE_PP0N_  clock_i _00392_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[266]\ _14393_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[253]$_DFFE_PP0N_  clock_i _00393_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[267]\ _14392_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[254]$_DFFE_PP0N_  clock_i _00394_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[268]\ _14391_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[255]$_DFFE_PP0N_  clock_i _00395_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[269]\ _14390_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[256]$_DFFE_PP0N_  clock_i _00396_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[270]\ _14389_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[257]$_DFFE_PP0N_  clock_i _00397_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[271]\ _14388_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[258]$_DFFE_PP0N_  clock_i _00398_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[6]\ _14387_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[259]$_DFFE_PP0N_  clock_i _00399_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[7]\ _14386_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[25]$_DFFE_PP0N_  clock_i _00400_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[7]\ _14385_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[260]$_DFFE_PP0N_  clock_i _00401_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[8]\ _14384_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[261]$_DFFE_PP0N_  clock_i _00402_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[9]\ _14383_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[262]$_DFFE_PP0N_  clock_i _00403_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[10]\ _14382_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[263]$_DFFE_PP0N_  clock_i _00404_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[11]\ _14381_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[264]$_DFFE_PP0N_  clock_i _00405_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[12]\ _14380_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[265]$_DFFE_PP0N_  clock_i _00406_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[13]\ _14379_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[266]$_DFFE_PP0N_  clock_i _00407_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[14]\ _14378_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[267]$_DFFE_PP0N_  clock_i _00408_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[15]\ _14377_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[268]$_DFFE_PP0N_  clock_i _00409_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[16]\ _14376_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[269]$_DFFE_PP0N_  clock_i _00410_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3008_o[17]\ _14375_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[26]$_DFFE_PP0N_  clock_i _00411_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[8]\ _14374_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[27]$_DFFE_PP0N_  clock_i _00412_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[9]\ _14373_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[28]$_DFFE_PP0N_  clock_i _00413_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[10]\ _14372_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[29]$_DFFE_PP0N_  clock_i _00414_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[11]\ _14371_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[2]$_DFFE_PP0N_  clock_i _00415_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[2]\ _14370_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[30]$_DFFE_PP0N_  clock_i _00416_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[12]\ _14369_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[31]$_DFFE_PP0N_  clock_i _00417_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[13]\ _14368_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[32]$_DFFE_PP0N_  clock_i _00418_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[14]\ _14367_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[33]$_DFFE_PP0N_  clock_i _00419_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[15]\ _14366_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[34]$_DFFE_PP0N_  clock_i _00420_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[16]\ _14365_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[35]$_DFFE_PP0N_  clock_i _00421_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2639_o[17]\ _14364_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[36]$_DFFE_PP0N_  clock_i _00422_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[38]\ _14363_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[37]$_DFFE_PP0N_  clock_i _00423_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[39]\ _14362_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[38]$_DFFE_PP0N_  clock_i _00424_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[40]\ _14361_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[39]$_DFFE_PP0N_  clock_i _00425_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[41]\ _14360_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[3]$_DFFE_PP0N_  clock_i _00426_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[3]\ _14359_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[40]$_DFFE_PP0N_  clock_i _00427_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[42]\ _14358_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[41]$_DFFE_PP0N_  clock_i _00428_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[43]\ _14357_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[42]$_DFFE_PP0N_  clock_i _00429_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[6]\ _14356_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[43]$_DFFE_PP0N_  clock_i _00430_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[7]\ _14355_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[44]$_DFFE_PP0N_  clock_i _00431_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[8]\ _14354_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[45]$_DFFE_PP0N_  clock_i _00432_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[9]\ _14353_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[46]$_DFFE_PP0N_  clock_i _00433_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[10]\ _14352_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[47]$_DFFE_PP0N_  clock_i _00434_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[11]\ _14351_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[48]$_DFFE_PP0N_  clock_i _00435_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[12]\ _14350_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[49]$_DFFE_PP0N_  clock_i _00436_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[13]\ _14349_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[4]$_DFFE_PP0N_  clock_i _00437_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[4]\ _14348_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[50]$_DFFE_PP0N_  clock_i _00438_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[14]\ _14347_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[51]$_DFFE_PP0N_  clock_i _00439_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[15]\ _14346_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[52]$_DFFE_PP0N_  clock_i _00440_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[16]\ _14345_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[53]$_DFFE_PP0N_  clock_i _00441_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2642_o[17]\ _14344_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[54]$_DFFE_PP0N_  clock_i _00442_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[57]\ _14343_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[55]$_DFFE_PP0N_  clock_i _00443_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[58]\ _14342_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[56]$_DFFE_PP0N_  clock_i _00444_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[59]\ _14341_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[57]$_DFFE_PP0N_  clock_i _00445_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[60]\ _14340_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[58]$_DFFE_PP0N_  clock_i _00446_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[61]\ _14339_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[59]$_DFFE_PP0N_  clock_i _00447_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[62]\ _14338_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[5]$_DFFE_PP0N_  clock_i _00448_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[5]\ _14337_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[60]$_DFFE_PP0N_  clock_i _00449_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[6]\ _14336_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[61]$_DFFE_PP0N_  clock_i _00450_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[7]\ _14335_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[62]$_DFFE_PP0N_  clock_i _00451_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[8]\ _14334_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[63]$_DFFE_PP0N_  clock_i _00452_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[9]\ _14333_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[64]$_DFFE_PP0N_  clock_i _00453_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[10]\ _14332_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[65]$_DFFE_PP0N_  clock_i _00454_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[11]\ _14331_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[66]$_DFFE_PP0N_  clock_i _00455_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[12]\ _14330_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[67]$_DFFE_PP0N_  clock_i _00456_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[13]\ _14329_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[68]$_DFFE_PP0N_  clock_i _00457_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[14]\ _14328_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[69]$_DFFE_PP0N_  clock_i _00458_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[15]\ _14327_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[6]$_DFFE_PP0N_  clock_i _00459_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[6]\ _14326_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[70]$_DFFE_PP0N_  clock_i _00460_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[16]\ _14325_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[71]$_DFFE_PP0N_  clock_i _00461_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2645_o[17]\ _14324_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[72]$_DFFE_PP0N_  clock_i _00462_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[76]\ _14323_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[73]$_DFFE_PP0N_  clock_i _00463_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[77]\ _14322_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[74]$_DFFE_PP0N_  clock_i _00464_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[78]\ _14321_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[75]$_DFFE_PP0N_  clock_i _00465_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[79]\ _14320_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[76]$_DFFE_PP0N_  clock_i _00466_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[80]\ _14319_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[77]$_DFFE_PP0N_  clock_i _00467_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[81]\ _14318_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[78]$_DFFE_PP0N_  clock_i _00468_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[6]\ _14317_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[79]$_DFFE_PP0N_  clock_i _00469_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[7]\ _14316_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[7]$_DFFE_PP0N_  clock_i _00470_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[7]\ _14315_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[80]$_DFFE_PP0N_  clock_i _00471_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[8]\ _14314_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[81]$_DFFE_PP0N_  clock_i _00472_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[9]\ _14313_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[82]$_DFFE_PP0N_  clock_i _00473_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[10]\ _14312_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[83]$_DFFE_PP0N_  clock_i _00474_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[11]\ _14311_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[84]$_DFFE_PP0N_  clock_i _00475_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[12]\ _14310_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[85]$_DFFE_PP0N_  clock_i _00476_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[13]\ _14309_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[86]$_DFFE_PP0N_  clock_i _00477_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[14]\ _14308_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[87]$_DFFE_PP0N_  clock_i _00478_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[15]\ _14307_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[88]$_DFFE_PP0N_  clock_i _00479_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[16]\ _14306_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[89]$_DFFE_PP0N_  clock_i _00480_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2648_o[17]\ _14305_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[8]$_DFFE_PP0N_  clock_i _00481_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[8]\ _14304_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[90]$_DFFE_PP0N_  clock_i _00482_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[95]\ _14303_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[91]$_DFFE_PP0N_  clock_i _00483_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[96]\ _14302_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[92]$_DFFE_PP0N_  clock_i _00484_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[97]\ _14301_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[93]$_DFFE_PP0N_  clock_i _00485_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[98]\ _14300_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[94]$_DFFE_PP0N_  clock_i _00486_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[99]\ _14299_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[95]$_DFFE_PP0N_  clock_i _00487_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.end_of_window_logic_virt_win_end[100]\ _14298_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[96]$_DFFE_PP0N_  clock_i _00488_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[6]\ _14297_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[97]$_DFFE_PP0N_  clock_i _00489_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[7]\ _14296_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[98]$_DFFE_PP0N_  clock_i _00490_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[8]\ _14295_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[99]$_DFFE_PP0N_  clock_i _00491_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2651_o[9]\ _14294_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3024_q[9]$_DFFE_PP0N_  clock_i _00492_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2636_o[9]\ _14293_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[0]$_DFFE_PP0P_  clock_i _00493_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2635_o[0]\ _00050_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[10]$_DFFE_PP0P_  clock_i _00494_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2650_o[0]\ _00041_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[11]$_DFFE_PP0P_  clock_i _00495_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2650_o[1]\ _14292_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[12]$_DFFE_PP0P_  clock_i _00496_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2653_o[0]\ _14291_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[13]$_DFFE_PP0P_  clock_i _00497_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2653_o[1]\ _14290_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[14]$_DFFE_PP0P_  clock_i _00498_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2656_o[0]\ _14289_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[15]$_DFFE_PP0P_  clock_i _00499_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2656_o[1]\ _14288_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[16]$_DFFE_PP0P_  clock_i _00500_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2659_o[0]\ _00106_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[17]$_DFFE_PP0P_  clock_i _00501_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2659_o[1]\ _14287_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[18]$_DFFE_PP0P_  clock_i _00502_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2662_o[0]\ _00105_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[19]$_DFFE_PP0P_  clock_i _00503_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2662_o[1]\ _14286_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[1]$_DFFE_PP0P_  clock_i _00504_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2635_o[1]\ _14285_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[20]$_DFFE_PP0P_  clock_i _00505_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2665_o[0]\ _00104_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[21]$_DFFE_PP0P_  clock_i _00506_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2665_o[1]\ _14284_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[22]$_DFFE_PP0P_  clock_i _00507_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2668_o[0]\ _00101_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[23]$_DFFE_PP0P_  clock_i _00508_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2668_o[1]\ _14283_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[24]$_DFFE_PP0P_  clock_i _00509_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2671_o[0]\ _00102_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[25]$_DFFE_PP0P_  clock_i _00510_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2671_o[1]\ _14282_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[26]$_DFFE_PP0P_  clock_i _00511_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2674_o[0]\ _00103_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[27]$_DFFE_PP0P_  clock_i _00512_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2674_o[1]\ _14281_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[28]$_DFFE_PP0P_  clock_i _00513_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n3499_o\ _14280_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[29]$_DFFE_PP0P_  clock_i _00514_ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.gen_spike_2_tc_n1_spike_2_tc.n3496_o\ _14279_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[2]$_DFFE_PP0P_  clock_i _00515_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2638_o[0]\ _00049_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[3]$_DFFE_PP0P_  clock_i _00516_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2638_o[1]\ _14278_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[4]$_DFFE_PP0P_  clock_i _00517_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2641_o[0]\ _00047_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[5]$_DFFE_PP0P_  clock_i _00518_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2641_o[1]\ _14277_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[6]$_DFFE_PP0P_  clock_i _00519_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2644_o[0]\ _00045_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[7]$_DFFE_PP0P_  clock_i _00520_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2644_o[1]\ _14276_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[8]$_DFFE_PP0P_  clock_i _00521_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2647_o[0]\ _00043_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3025_q[9]$_DFFE_PP0P_  clock_i _00522_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2647_o[1]\ _14275_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[0]$_DFFE_PP0P_  clock_i _00523_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2637_o\ _14274_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[10]$_DFFE_PP0P_  clock_i _00524_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2667_o\ _14273_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[11]$_DFFE_PP0P_  clock_i _00525_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2670_o\ _14272_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[12]$_DFFE_PP0P_  clock_i _00526_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2673_o\ _14271_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[13]$_DFFE_PP0P_  clock_i _00527_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2676_o\ _14270_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[14]$_DFFE_PP0P_  clock_i _00528_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3011_o\ _14269_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[1]$_DFFE_PP0P_  clock_i _00529_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2640_o\ _14268_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[2]$_DFFE_PP0P_  clock_i _00530_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2643_o\ _14267_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[3]$_DFFE_PP0P_  clock_i _00531_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2646_o\ _14266_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[4]$_DFFE_PP0P_  clock_i _00532_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2649_o\ _14265_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[5]$_DFFE_PP0P_  clock_i _00533_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2652_o\ _14264_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[6]$_DFFE_PP0P_  clock_i _00534_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2655_o\ _14263_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[7]$_DFFE_PP0P_  clock_i _00535_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2658_o\ _14262_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[8]$_DFFE_PP0P_  clock_i _00536_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2661_o\ _14261_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3027_q[9]$_DFFE_PP0P_  clock_i _00537_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2664_o\ _14260_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3028_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n2778_o\ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.n3028_q\ _14259_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[48]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[0]\ _00040_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[49]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[1]\ _00042_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[2]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[50]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[2]\ _00044_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[3]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[51]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[3]\ _00046_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[4]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[52]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[4]\ _00048_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3236_q[5]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_thermocodes[53]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.buf_reg[5]\ _14258_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3237_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.n1658_o\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3033_o\ _14257_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3237_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3033_o\ \atbs_core_0.adaptive_ctrl_0.n1689_o\ _14256_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[0]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[0]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[0]\ _14255_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[1]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[1]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[1]\ _14254_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[2]$_DFF_PP0_  clock_i \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3234_o[2]\ \atbs_core_0.adaptive_ctrl_0.weyls_discrepancy_0.n3242_q[2]\ _14253_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[0]$_DFFE_PP0P_  clock_i _00538_ \atbs_core_0.analog_trigger_0.counter_value[0]\ _14252_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[1]$_DFFE_PP0P_  clock_i _00539_ \atbs_core_0.analog_trigger_0.counter_value[1]\ _14251_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[2]$_DFFE_PP0P_  clock_i _00540_ \atbs_core_0.analog_trigger_0.counter_value[2]\ _14250_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[3]$_DFFE_PP0P_  clock_i _00541_ \atbs_core_0.analog_trigger_0.counter_value[3]\ _14249_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[4]$_DFFE_PP0P_  clock_i _00542_ \atbs_core_0.analog_trigger_0.counter_value[4]\ _14248_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[5]$_DFFE_PP0P_  clock_i _00543_ \atbs_core_0.analog_trigger_0.counter_value[5]\ _14247_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.analog_trigger_0.n2120_q[6]$_DFFE_PP0P_  clock_i _00544_ \atbs_core_0.analog_trigger_0.counter_value[6]\ _14246_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1937_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1836_o\ \atbs_core_0.dac_control_0.n1833_o\ _14245_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1938_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1833_o\ \atbs_core_0.dac_control_0.n1938_q\ _00094_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[1]$_DFFE_PP0N_  clock_i _00545_ \atbs_core_0.dac_control_0.dac_init_value[1]\ _14244_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[2]$_DFFE_PP0N_  clock_i _00546_ \atbs_core_0.dac_control_0.dac_init_value[2]\ _14243_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[3]$_DFFE_PP0N_  clock_i _00547_ \atbs_core_0.dac_control_0.dac_init_value[3]\ _14242_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[4]$_DFFE_PP0N_  clock_i _00548_ \atbs_core_0.dac_control_0.dac_init_value[4]\ _14241_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[5]$_DFFE_PP0N_  clock_i _00549_ \atbs_core_0.dac_control_0.dac_init_value[5]\ _14240_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[6]$_DFFE_PP0N_  clock_i _00550_ \atbs_core_0.dac_control_0.dac_init_value[6]\ _14239_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1939_q[7]$_DFFE_PP0N_  clock_i _00551_ \atbs_core_0.dac_control_0.dac_init_value[7]\ _14238_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[0]$_DFFE_PP0P_  clock_i _00552_ \atbs_core_0.dac_control_0.dac_counter_value[0]\ _00037_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[1]$_DFFE_PP0P_  clock_i _00553_ \atbs_core_0.dac_control_0.dac_counter_value[1]\ _00079_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[2]$_DFFE_PP0P_  clock_i _00554_ \atbs_core_0.dac_control_0.dac_counter_value[2]\ _00083_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[3]$_DFFE_PP0P_  clock_i _00555_ \atbs_core_0.dac_control_0.dac_counter_value[3]\ _00089_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[4]$_DFFE_PP0P_  clock_i _00556_ \atbs_core_0.dac_control_0.dac_counter_value[4]\ _00087_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[5]$_DFFE_PP0P_  clock_i _00557_ \atbs_core_0.dac_control_0.dac_counter_value[5]\ _00085_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[6]$_DFFE_PP0P_  clock_i _00558_ \atbs_core_0.dac_control_0.dac_counter_value[6]\ _00038_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1940_q[7]$_DFFE_PP0P_  clock_i _00559_ \atbs_core_0.dac_control_0.dac_counter_value[7]\ _00093_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1941_q$_DFFE_PP0P_  clock_i _00560_ \atbs_core_0.dac_control_0.dac_change_in_progress\ _14237_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1942_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1904_o[0]\ \atbs_core_0.dac_control_0.n1942_q[0]\ _14236_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1942_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1904_o[1]\ \atbs_core_0.dac_control_0.n1942_q[1]\ _14235_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1942_q[2]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.n1904_o[2]\ \atbs_core_0.dac_control_0.n1942_q[2]\ _00058_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1943_q[0]$_DFFE_PP0P_  clock_i _00561_ dac_upper_o[0] _14234_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1943_q[1]$_DFFE_PP0P_  clock_i _00562_ dac_upper_o[1] _14233_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1943_q[2]$_DFFE_PP0P_  clock_i _00563_ dac_upper_o[2] _14232_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.n1943_q[3]$_DFFE_PP0P_  clock_i _00564_ dac_upper_o[3] _14231_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.sync_chain_0.async_i\ \atbs_core_0.dac_control_0.sync_chain_0.n1426_o\ _14230_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_0.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_0.sync_chain_0.n1426_o\ \atbs_core_0.dac_control_0.n1913_o\ _14229_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2086_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1984_o\ \atbs_core_0.dac_control_1.n1981_o\ _14228_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2087_q$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n1981_o\ \atbs_core_0.dac_control_1.n2087_q\ _00099_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2088_q[6]$_DFFE_PP0N_  clock_i _00565_ \atbs_core_0.dac_control_1.dac_init_value[6]\ _14227_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[0]$_DFFE_PP0P_  clock_i _00566_ \atbs_core_0.dac_control_1.dac_counter_value[0]\ _14226_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[1]$_DFFE_PP0P_  clock_i _00567_ \atbs_core_0.dac_control_1.dac_counter_value[1]\ _00097_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[2]$_DFFE_PP0P_  clock_i _00568_ \atbs_core_0.dac_control_1.dac_counter_value[2]\ _00096_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[3]$_DFFE_PP0P_  clock_i _00569_ \atbs_core_0.dac_control_1.dac_counter_value[3]\ _00095_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[4]$_DFFE_PP0P_  clock_i _00570_ \atbs_core_0.dac_control_1.dac_counter_value[4]\ _00098_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[5]$_DFFE_PP0P_  clock_i _00571_ \atbs_core_0.dac_control_1.dac_counter_value[5]\ _14225_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[6]$_DFFE_PP0P_  clock_i _00572_ \atbs_core_0.dac_control_1.dac_counter_value[6]\ _14224_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2089_q[7]$_DFFE_PP0P_  clock_i _00573_ \atbs_core_0.dac_control_1.dac_counter_value[7]\ _00036_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2090_q$_DFFE_PP0P_  clock_i _00574_ \atbs_core_0.dac_control_1.dac_change_in_progress\ _14223_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2091_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n2053_o[0]\ \atbs_core_0.dac_control_1.n2091_q[0]\ _14222_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2091_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n2053_o[1]\ \atbs_core_0.dac_control_1.n2091_q[1]\ _14221_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2091_q[2]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.n2053_o[2]\ \atbs_core_0.dac_control_1.n2091_q[2]\ _00059_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2092_q[0]$_DFFE_PP0P_  clock_i _00575_ dac_lower_o[0] _14220_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2092_q[1]$_DFFE_PP0P_  clock_i _00576_ dac_lower_o[1] _14219_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2092_q[2]$_DFFE_PP0P_  clock_i _00577_ dac_lower_o[2] _14218_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.n2092_q[3]$_DFFE_PP0P_  clock_i _00578_ dac_lower_o[3] _14217_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.sync_chain_0.async_i\ \atbs_core_0.dac_control_1.sync_chain_0.n1426_o\ _14216_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.dac_control_1.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.dac_control_1.sync_chain_0.n1426_o\ \atbs_core_0.dac_control_1.n2062_o\ _14215_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.bouncing_sync\ \atbs_core_0.debouncer_0.bouncing_sync_d\ _14214_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[0]\ \atbs_core_0.debouncer_0.counter_value[0]\ _14213_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[10]\ \atbs_core_0.debouncer_0.counter_value[10]\ _14212_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[11]\ \atbs_core_0.debouncer_0.counter_value[11]\ _14211_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[12]\ \atbs_core_0.debouncer_0.counter_value[12]\ _14210_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[13]\ \atbs_core_0.debouncer_0.counter_value[13]\ _14209_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[14]\ \atbs_core_0.debouncer_0.counter_value[14]\ _14208_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[15]\ \atbs_core_0.debouncer_0.counter_value[15]\ _14207_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[1]\ \atbs_core_0.debouncer_0.counter_value[1]\ _14206_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[2]\ \atbs_core_0.debouncer_0.counter_value[2]\ _14205_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[3]\ \atbs_core_0.debouncer_0.counter_value[3]\ _14204_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[4]\ \atbs_core_0.debouncer_0.counter_value[4]\ _14203_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[5]\ \atbs_core_0.debouncer_0.counter_value[5]\ _14202_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[6]\ \atbs_core_0.debouncer_0.counter_value[6]\ _14201_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[7]\ \atbs_core_0.debouncer_0.counter_value[7]\ _14200_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[8]\ \atbs_core_0.debouncer_0.counter_value[8]\ _14199_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.n1466_o[9]\ \atbs_core_0.debouncer_0.counter_value[9]\ _14198_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1511_q[0]$_DFFE_PP0P_  clock_i _00579_ \atbs_core_0.debouncer_0.n1511_q[0]\ _14197_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1511_q[1]$_DFFE_PP0P_  clock_i _00580_ \atbs_core_0.debouncer_0.n1511_q[1]\ _14196_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.n1512_q$_DFFE_PP0P_  clock_i _00581_ \atbs_core_0.debouncer_0.debounced\ _14195_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i trigger_start_mode_i \atbs_core_0.debouncer_0.sync_chain_0.n1426_o\ _14194_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_0.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_0.bouncing_sync\ _14193_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.bouncing_sync\ \atbs_core_0.debouncer_1.bouncing_sync_d\ _14192_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[0]\ \atbs_core_0.debouncer_1.counter_value[0]\ _14191_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[10]\ \atbs_core_0.debouncer_1.counter_value[10]\ _14190_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[11]\ \atbs_core_0.debouncer_1.counter_value[11]\ _14189_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[12]\ \atbs_core_0.debouncer_1.counter_value[12]\ _14188_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[13]\ \atbs_core_0.debouncer_1.counter_value[13]\ _14187_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[14]\ \atbs_core_0.debouncer_1.counter_value[14]\ _14186_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[15]\ \atbs_core_0.debouncer_1.counter_value[15]\ _14185_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[1]\ \atbs_core_0.debouncer_1.counter_value[1]\ _14184_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[2]\ \atbs_core_0.debouncer_1.counter_value[2]\ _14183_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[3]\ \atbs_core_0.debouncer_1.counter_value[3]\ _14182_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[4]\ \atbs_core_0.debouncer_1.counter_value[4]\ _14181_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[5]\ \atbs_core_0.debouncer_1.counter_value[5]\ _14180_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[6]\ \atbs_core_0.debouncer_1.counter_value[6]\ _14179_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[7]\ \atbs_core_0.debouncer_1.counter_value[7]\ _14178_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[8]\ \atbs_core_0.debouncer_1.counter_value[8]\ _14177_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.n1466_o[9]\ \atbs_core_0.debouncer_1.counter_value[9]\ _14176_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1511_q[0]$_DFFE_PP0P_  clock_i _00582_ \atbs_core_0.debouncer_1.n1511_q[0]\ _14175_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1511_q[1]$_DFFE_PP0P_  clock_i _00583_ \atbs_core_0.debouncer_1.n1511_q[1]\ _14174_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.n1512_q$_DFFE_PP0P_  clock_i _00584_ \atbs_core_0.adaptive_mode_debounced\ _14173_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i adaptive_mode_i \atbs_core_0.debouncer_1.sync_chain_0.n1426_o\ _14172_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_1.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_1.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_1.bouncing_sync\ _14171_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.bouncing_sync\ \atbs_core_0.debouncer_2.bouncing_sync_d\ _14170_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[0]\ \atbs_core_0.debouncer_2.counter_value[0]\ _14169_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[10]\ \atbs_core_0.debouncer_2.counter_value[10]\ _14168_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[11]\ \atbs_core_0.debouncer_2.counter_value[11]\ _14167_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[12]\ \atbs_core_0.debouncer_2.counter_value[12]\ _14166_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[13]\ \atbs_core_0.debouncer_2.counter_value[13]\ _14165_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[14]\ \atbs_core_0.debouncer_2.counter_value[14]\ _14164_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[15]\ \atbs_core_0.debouncer_2.counter_value[15]\ _14163_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[1]\ \atbs_core_0.debouncer_2.counter_value[1]\ _14162_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[2]\ \atbs_core_0.debouncer_2.counter_value[2]\ _14161_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[3]\ \atbs_core_0.debouncer_2.counter_value[3]\ _14160_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[4]\ \atbs_core_0.debouncer_2.counter_value[4]\ _14159_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[5]\ \atbs_core_0.debouncer_2.counter_value[5]\ _14158_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[6]\ \atbs_core_0.debouncer_2.counter_value[6]\ _14157_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[7]\ \atbs_core_0.debouncer_2.counter_value[7]\ _14156_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[8]\ \atbs_core_0.debouncer_2.counter_value[8]\ _14155_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.n1466_o[9]\ \atbs_core_0.debouncer_2.counter_value[9]\ _14154_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1511_q[0]$_DFFE_PP0P_  clock_i _00585_ \atbs_core_0.debouncer_2.n1511_q[0]\ _14153_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1511_q[1]$_DFFE_PP0P_  clock_i _00586_ \atbs_core_0.debouncer_2.n1511_q[1]\ _14152_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.n1512_q$_DFFE_PP0P_  clock_i _00587_ \atbs_core_0.control_mode_debounced\ _14151_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i control_mode_i \atbs_core_0.debouncer_2.sync_chain_0.n1426_o\ _14150_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_2.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_2.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_2.bouncing_sync\ _14149_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.bouncing_sync\ \atbs_core_0.debouncer_3.bouncing_sync_d\ _14148_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[0]\ \atbs_core_0.debouncer_3.counter_value[0]\ _14147_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[10]\ \atbs_core_0.debouncer_3.counter_value[10]\ _14146_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[11]\ \atbs_core_0.debouncer_3.counter_value[11]\ _14145_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[12]\ \atbs_core_0.debouncer_3.counter_value[12]\ _14144_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[13]\ \atbs_core_0.debouncer_3.counter_value[13]\ _14143_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[14]\ \atbs_core_0.debouncer_3.counter_value[14]\ _14142_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[15]\ \atbs_core_0.debouncer_3.counter_value[15]\ _14141_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[1]\ \atbs_core_0.debouncer_3.counter_value[1]\ _14140_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[2]\ \atbs_core_0.debouncer_3.counter_value[2]\ _14139_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[3]\ \atbs_core_0.debouncer_3.counter_value[3]\ _14138_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[4]\ \atbs_core_0.debouncer_3.counter_value[4]\ _14137_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[5]\ \atbs_core_0.debouncer_3.counter_value[5]\ _14136_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[6]\ \atbs_core_0.debouncer_3.counter_value[6]\ _14135_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[7]\ \atbs_core_0.debouncer_3.counter_value[7]\ _14134_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[8]\ \atbs_core_0.debouncer_3.counter_value[8]\ _14133_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.n1466_o[9]\ \atbs_core_0.debouncer_3.counter_value[9]\ _14132_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1511_q[0]$_DFFE_PP0P_  clock_i _00588_ \atbs_core_0.debouncer_3.n1511_q[0]\ _14131_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1511_q[1]$_DFFE_PP0P_  clock_i _00589_ \atbs_core_0.debouncer_3.n1511_q[1]\ _14130_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.n1512_q$_DFFE_PP0P_  clock_i _00590_ \atbs_core_0.debouncer_3.debounced\ _00039_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i signal_select_in_i \atbs_core_0.debouncer_3.sync_chain_0.n1426_o\ _14129_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_3.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_3.bouncing_sync\ _14128_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.bouncing_sync\ \atbs_core_0.debouncer_4.bouncing_sync_d\ _14127_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[0]\ \atbs_core_0.debouncer_4.counter_value[0]\ _14126_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[10]\ \atbs_core_0.debouncer_4.counter_value[10]\ _14125_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[11]\ \atbs_core_0.debouncer_4.counter_value[11]\ _14124_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[12]\ \atbs_core_0.debouncer_4.counter_value[12]\ _14123_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[13]\ \atbs_core_0.debouncer_4.counter_value[13]\ _14122_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[14]\ \atbs_core_0.debouncer_4.counter_value[14]\ _14121_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[15]\ \atbs_core_0.debouncer_4.counter_value[15]\ _14120_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[1]\ \atbs_core_0.debouncer_4.counter_value[1]\ _14119_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[2]\ \atbs_core_0.debouncer_4.counter_value[2]\ _14118_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[3]\ \atbs_core_0.debouncer_4.counter_value[3]\ _14117_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[4]\ \atbs_core_0.debouncer_4.counter_value[4]\ _14116_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[5]\ \atbs_core_0.debouncer_4.counter_value[5]\ _14115_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[6]\ \atbs_core_0.debouncer_4.counter_value[6]\ _14114_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[7]\ \atbs_core_0.debouncer_4.counter_value[7]\ _14113_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[8]\ \atbs_core_0.debouncer_4.counter_value[8]\ _14112_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.n1466_o[9]\ \atbs_core_0.debouncer_4.counter_value[9]\ _14111_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1511_q[0]$_DFFE_PP0P_  clock_i _00591_ \atbs_core_0.debouncer_4.n1511_q[0]\ _14110_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1511_q[1]$_DFFE_PP0P_  clock_i _00592_ \atbs_core_0.debouncer_4.n1511_q[1]\ _14109_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.n1512_q$_DFFE_PP0P_  clock_i _00593_ \atbs_core_0.debouncer_4.debounced\ _14108_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i enable_i \atbs_core_0.debouncer_4.sync_chain_0.n1426_o\ _14107_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_4.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_4.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_4.bouncing_sync\ _14106_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1509_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.bouncing_sync\ \atbs_core_0.debouncer_5.bouncing_sync_d\ _14105_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[0]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[0]\ \atbs_core_0.debouncer_5.counter_value[0]\ _14104_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[10]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[10]\ \atbs_core_0.debouncer_5.counter_value[10]\ _14103_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[11]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[11]\ \atbs_core_0.debouncer_5.counter_value[11]\ _14102_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[12]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[12]\ \atbs_core_0.debouncer_5.counter_value[12]\ _14101_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[13]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[13]\ \atbs_core_0.debouncer_5.counter_value[13]\ _14100_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[14]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[14]\ \atbs_core_0.debouncer_5.counter_value[14]\ _14099_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[15]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[15]\ \atbs_core_0.debouncer_5.counter_value[15]\ _14098_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[1]\ \atbs_core_0.debouncer_5.counter_value[1]\ _14097_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[2]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[2]\ \atbs_core_0.debouncer_5.counter_value[2]\ _14096_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[3]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[3]\ \atbs_core_0.debouncer_5.counter_value[3]\ _14095_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[4]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[4]\ \atbs_core_0.debouncer_5.counter_value[4]\ _14094_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[5]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[5]\ \atbs_core_0.debouncer_5.counter_value[5]\ _14093_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[6]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[6]\ \atbs_core_0.debouncer_5.counter_value[6]\ _14092_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[7]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[7]\ \atbs_core_0.debouncer_5.counter_value[7]\ _14091_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[8]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[8]\ \atbs_core_0.debouncer_5.counter_value[8]\ _14090_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1510_q[9]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.n1466_o[9]\ \atbs_core_0.debouncer_5.counter_value[9]\ _14089_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1511_q[0]$_DFFE_PP0P_  clock_i _00594_ \atbs_core_0.debouncer_5.n1511_q[0]\ _14088_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1511_q[1]$_DFFE_PP0P_  clock_i _00595_ \atbs_core_0.debouncer_5.n1511_q[1]\ _14087_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.n1512_q$_DFFE_PP0P_  clock_i _00596_ \atbs_core_0.debouncer_5.debounced\ _14086_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.sync_chain_0.n1433_q[0]$_DFF_PP0_  clock_i select_tbs_delta_steps_i \atbs_core_0.debouncer_5.sync_chain_0.n1426_o\ _14085_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.debouncer_5.sync_chain_0.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.sync_chain_0.n1426_o\ \atbs_core_0.debouncer_5.bouncing_sync\ _14084_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[0]$_DFFE_PP0P_  clock_i _00597_ \atbs_core_0.uart_0.uart_tx_0.n3348_o\ _14083_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[10]$_DFFE_PP0P_  clock_i _00598_ \atbs_core_0.memory2uart_0.n2574_o[2]\ _14082_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[11]$_DFFE_PP0P_  clock_i _00599_ \atbs_core_0.memory2uart_0.n2574_o[3]\ _14081_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[12]$_DFFE_PP0P_  clock_i _00600_ \atbs_core_0.memory2uart_0.n2574_o[4]\ _14080_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[13]$_DFFE_PP0P_  clock_i _00601_ \atbs_core_0.memory2uart_0.n2574_o[5]\ _14079_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[14]$_DFFE_PP0P_  clock_i _00602_ \atbs_core_0.memory2uart_0.n2574_o[6]\ _14078_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[15]$_DFFE_PP0P_  clock_i _00603_ \atbs_core_0.memory2uart_0.n2574_o[7]\ _14077_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[16]$_DFFE_PP0P_  clock_i _00604_ \atbs_core_0.memory2uart_0.n2574_o[8]\ _14076_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[17]$_DFFE_PP0P_  clock_i _00605_ \atbs_core_0.memory2uart_0.n2574_o[9]\ _14075_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[18]$_DFFE_PP0P_  clock_i _00606_ \atbs_core_0.memory2uart_0.n2574_o[10]\ _14074_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[19]$_DFFE_PP0P_  clock_i _00607_ \atbs_core_0.memory2uart_0.n2574_o[11]\ _14073_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[1]$_DFFE_PP0P_  clock_i _00608_ \atbs_core_0.uart_0.uart_tx_0.n3349_o\ _14072_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[20]$_DFFE_PP0P_  clock_i _00609_ \atbs_core_0.memory2uart_0.n2574_o[12]\ _14071_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[21]$_DFFE_PP0P_  clock_i _00610_ \atbs_core_0.memory2uart_0.n2574_o[13]\ _14070_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[22]$_DFFE_PP0P_  clock_i _00611_ \atbs_core_0.memory2uart_0.n2574_o[14]\ _14069_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[23]$_DFFE_PP0P_  clock_i _00612_ \atbs_core_0.memory2uart_0.n2574_o[15]\ _14068_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[2]$_DFFE_PP0P_  clock_i _00613_ \atbs_core_0.uart_0.uart_tx_0.n3350_o\ _14067_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[3]$_DFFE_PP0P_  clock_i _00614_ \atbs_core_0.uart_0.uart_tx_0.n3351_o\ _14066_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[4]$_DFFE_PP0P_  clock_i _00615_ \atbs_core_0.uart_0.uart_tx_0.n3352_o\ _14065_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[5]$_DFFE_PP0P_  clock_i _00616_ \atbs_core_0.uart_0.uart_tx_0.n3353_o\ _14064_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[6]$_DFFE_PP0P_  clock_i _00617_ \atbs_core_0.uart_0.uart_tx_0.n3354_o\ _14063_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[7]$_DFFE_PP0P_  clock_i _00618_ \atbs_core_0.uart_0.uart_tx_0.n3355_o\ _14062_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[8]$_DFFE_PP0P_  clock_i _00619_ \atbs_core_0.memory2uart_0.n2574_o[0]\ _14061_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2603_q[9]$_DFFE_PP0P_  clock_i _00620_ \atbs_core_0.memory2uart_0.n2574_o[1]\ _14060_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2605_q$_DFF_PP0_  clock_i \atbs_core_0.memory2uart_0.n2588_o\ \atbs_core_0.memory2uart_0.n2605_q\ _00062_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2606_q[0]$_DFFE_PP0P_  clock_i _00621_ \atbs_core_0.memory2uart_0.counter[0]\ _14059_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.memory2uart_0.n2606_q[1]$_DFFE_PP0P_  clock_i _00622_ \atbs_core_0.memory2uart_0.counter[1]\ _14058_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1379_q$_DFF_PP0_  clock_i \atbs_core_0.adaptive_mode_debounced\ \atbs_core_0.adaptive_mode_d\ _14057_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1380_q$_DFF_PP0_  clock_i \atbs_core_0.control_mode_debounced\ \atbs_core_0.control_mode_d\ _14056_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1381_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_3.debounced\ \atbs_core_0.n1381_q\ _14055_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1382_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_5.debounced\ \atbs_core_0.n1382_q\ _14054_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1383_q$_DFF_PP0_  clock_i \atbs_core_0.debouncer_0.debounced\ \atbs_core_0.n1383_q\ _14053_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1384_q$_DFF_PP0_  clock_i \atbs_core_0.n72_o\ \atbs_core_0.n1384_q\ _14052_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1385_q$_DFFE_PP0P_  clock_i _00623_ \atbs_core_0.detection_en\ _14051_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1386_q$_DFF_PP0_  clock_i \atbs_core_0.n179_o\ \atbs_core_0.n1386_q\ _14050_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1387_q$_DFF_PP0_  clock_i \atbs_core_0.n187_o\ \atbs_core_0.n1387_q\ _14049_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1388_q$_DFFE_PP0P_  clock_i _00624_ \atbs_core_0.clear_dac\ _14048_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1389_q$_DFFE_PP0P_  clock_i _00625_ \atbs_core_0.n1389_q\ _14047_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1390_q$_DFFE_PP0P_  clock_i _00626_ \atbs_core_0.enable_read\ _14046_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1391_q$_DFFE_PP0P_  clock_i _00627_ \atbs_core_0.analog_trigger_uart\ _14045_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1392_q[3]$_DFFE_PP0P_  clock_i _00628_ \atbs_core_0.analog_trigger_0.period_adj_i[3]\ _14044_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1392_q[4]$_DFFE_PP0P_  clock_i _00629_ \atbs_core_0.analog_trigger_0.period_adj_i[4]\ _14043_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1392_q[5]$_DFFE_PP0P_  clock_i _00630_ \atbs_core_0.analog_trigger_0.period_adj_i[5]\ _14042_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1392_q[6]$_DFFE_PP0P_  clock_i _00631_ \atbs_core_0.analog_trigger_0.period_adj_i[6]\ _14041_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1393_q$_DFFE_PP0P_  clock_i _00632_ \atbs_core_0.n1393_q\ _00060_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1394_q[6]$_DFFE_PP1P_  clock_i _00633_ _00164_ \atbs_core_0.n1394_q[6]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1394_q[7]$_DFFE_PP0P_  clock_i _00634_ \atbs_core_0.n1394_q[7]\ _14040_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1395_q$_DFFE_PP0P_  clock_i _00635_ \atbs_core_0.n1395_q\ _14039_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1396_q[6]$_DFFE_PP1P_  clock_i _00636_ _00165_ \atbs_core_0.n1396_q[6]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1396_q[7]$_DFFE_PP0P_  clock_i _00637_ \atbs_core_0.n1396_q[7]\ _14038_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1397_q$_DFFE_PP0P_  clock_i _00638_ \atbs_core_0.n1397_q\ _00066_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1398_q[6]$_DFFE_PP1P_  clock_i _00639_ _00166_ \atbs_core_0.n1398_q[6]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1398_q[7]$_DFFE_PP0P_  clock_i _00640_ \atbs_core_0.n1398_q[7]\ _14037_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1399_q$_DFFE_PP0P_  clock_i _00641_ \atbs_core_0.n1399_q\ _14036_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1400_q[10]$_DFFE_PP0P_  clock_i _00642_ \atbs_core_0.n1400_q[10]\ _14035_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1401_q$_DFFE_PP0P_  clock_i _00643_ \atbs_core_0.n1401_q\ _00107_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1402_q[0]$_DFFE_PP1P_  clock_i _00644_ _00167_ \atbs_core_0.n1402_q[0]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1402_q[1]$_DFFE_PP1P_  clock_i _00645_ _00168_ \atbs_core_0.n1402_q[1]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1402_q[2]$_DFFE_PP1P_  clock_i _00646_ _00169_ \atbs_core_0.n1402_q[2]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1403_q$_DFFE_PP0P_  clock_i _00647_ \atbs_core_0.baudrate_uart\ _00064_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[0]$_DFFE_PP1P_  clock_i _00648_ _00170_ \atbs_core_0.baudrate_adj_uart[0]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[2]$_DFFE_PP1P_  clock_i _00649_ _00171_ \atbs_core_0.baudrate_adj_uart[2]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[3]$_DFFE_PP0P_  clock_i _00650_ \atbs_core_0.baudrate_adj_uart[1]\ _14034_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[4]$_DFFE_PP0P_  clock_i _00651_ \atbs_core_0.baudrate_adj_uart[4]\ _14033_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[5]$_DFFE_PP0P_  clock_i _00652_ \atbs_core_0.baudrate_adj_uart[5]\ _14032_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[6]$_DFFE_PP1P_  clock_i _00653_ _00172_ \atbs_core_0.baudrate_adj_uart[6]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1404_q[7]$_DFFE_PP0P_  clock_i _00654_ \atbs_core_0.baudrate_adj_uart[7]\ _14031_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1405_q$_DFFE_PP0P_  clock_i _00655_ \atbs_core_0.n1405_q\ _00065_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1406_q[1]$_DFFE_PP0P_  clock_i _00656_ \atbs_core_0.n1406_q[1]\ _14030_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1406_q[2]$_DFFE_PP1P_  clock_i _00657_ _00173_ \atbs_core_0.n1406_q[2]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1406_q[3]$_DFFE_PP0P_  clock_i _00658_ \atbs_core_0.n1406_q[3]\ _14029_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1406_q[4]$_DFFE_PP0P_  clock_i _00659_ \atbs_core_0.n1406_q[4]\ _14028_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1407_q$_DFFE_PP0P_  clock_i _00660_ \atbs_core_0.atbs_win_length_uart\ _14027_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[10]$_DFFE_PP1P_  clock_i _00661_ _00174_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[10]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[11]$_DFFE_PP1P_  clock_i _00662_ _00175_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[11]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[12]$_DFFE_PP1P_  clock_i _00663_ _00176_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[12]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[13]$_DFFE_PP1P_  clock_i _00664_ _00177_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[13]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[14]$_DFFE_PP1P_  clock_i _00665_ _00178_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[14]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[15]$_DFFE_PP0P_  clock_i _00666_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[15]\ _14026_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[16]$_DFFE_PP0P_  clock_i _00667_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[16]\ _14025_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[17]$_DFFE_PP0P_  clock_i _00668_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[17]\ _14024_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[6]$_DFFE_PP0P_  clock_i _00669_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[6]\ _14023_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[7]$_DFFE_PP0P_  clock_i _00670_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[7]\ _14022_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[8]$_DFFE_PP1P_  clock_i _00671_ _00179_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[8]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1408_q[9]$_DFFE_PP0P_  clock_i _00672_ \atbs_core_0.adaptive_ctrl_0.spike_shift_reg_0.win_length_i[9]\ _14021_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1409_q$_DFFE_PP0P_  clock_i _00673_ \atbs_core_0.atbs_max_delta_steps_uart\ _00108_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1410_q[1]$_DFFE_PP0P_  clock_i _00674_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[1]\ _14020_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1410_q[2]$_DFFE_PP0P_  clock_i _00675_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[2]\ _14019_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1410_q[3]$_DFFE_PP0P_  clock_i _00676_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[3]\ _14018_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1410_q[4]$_DFFE_PP1P_  clock_i _00677_ _00180_ \atbs_core_0.adaptive_ctrl_0.max_delta_steps_i[4]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[0]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[0]\ \atbs_core_0.main_counter_value[0]\ _14017_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[10]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[10]\ \atbs_core_0.main_counter_value[10]\ _14016_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[11]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[11]\ \atbs_core_0.main_counter_value[11]\ _14015_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[12]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[12]\ \atbs_core_0.main_counter_value[12]\ _14014_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[13]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[13]\ \atbs_core_0.main_counter_value[13]\ _14013_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[14]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[14]\ \atbs_core_0.main_counter_value[14]\ _14012_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[15]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[15]\ \atbs_core_0.main_counter_value[15]\ _14011_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[16]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[16]\ \atbs_core_0.main_counter_value[16]\ _14010_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[17]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[17]\ \atbs_core_0.main_counter_value[17]\ _14009_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[18]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[18]\ \atbs_core_0.main_counter_value[18]\ _14008_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[19]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[19]\ \atbs_core_0.main_counter_value[19]\ _14007_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[1]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[1]\ \atbs_core_0.main_counter_value[1]\ _14006_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[2]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[2]\ \atbs_core_0.main_counter_value[2]\ _14005_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[3]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[3]\ \atbs_core_0.main_counter_value[3]\ _14004_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[4]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[4]\ \atbs_core_0.main_counter_value[4]\ _14003_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[5]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[5]\ \atbs_core_0.main_counter_value[5]\ _14002_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[6]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[6]\ \atbs_core_0.main_counter_value[6]\ _14001_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[7]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[7]\ \atbs_core_0.main_counter_value[7]\ _14000_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[8]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[8]\ \atbs_core_0.main_counter_value[8]\ _13999_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1411_q[9]$_DFF_PP0_  clock_i \atbs_core_0.n268_o[9]\ \atbs_core_0.main_counter_value[9]\ _13998_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1412_q[0]$_DFF_PP1_  clock_i _00187_ _14574_ \atbs_core_0.n1412_q[0]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1412_q[1]$_DFF_PP0_  clock_i \atbs_core_0.n453_o[1]\ \atbs_core_0.n1412_q[1]\ _13997_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1412_q[2]$_DFF_PP0_  clock_i \atbs_core_0.n453_o[2]\ \atbs_core_0.n1412_q[2]\ _00056_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1413_q$_DFFE_PP0P_  clock_i _00678_ idle_led_o _13996_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1414_q$_DFFE_PP0P_  clock_i _00679_ overflow_led_o _13995_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1415_q$_DFFE_PP0P_  clock_i _00680_ underflow_led_o _13994_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1416_q$_DFFE_PP1P_  clock_i _00681_ _00181_ \atbs_core_0.n1416_q\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1417_q$_DFFE_PP0P_  clock_i _00682_ \atbs_core_0.adaptive_mode_uart\ _13993_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1418_q$_DFFE_PP1P_  clock_i _00683_ _00182_ \atbs_core_0.n1418_q\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1419_q$_DFFE_PP1P_  clock_i _00684_ _00183_ \atbs_core_0.enable_analog_uart\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.n1420_q$_DFFE_PP1P_  clock_i _00685_ _00184_ \atbs_core_0.n1420_q\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[0]$_DFFE_PP0P_  clock_i _00686_ \atbs_core_0.sc_noc_generator_0.counter_value[0]\ _13992_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[1]$_DFFE_PP0P_  clock_i _00687_ \atbs_core_0.sc_noc_generator_0.counter_value[1]\ _13991_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[2]$_DFFE_PP0P_  clock_i _00688_ \atbs_core_0.sc_noc_generator_0.counter_value[2]\ _13990_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[3]$_DFFE_PP0P_  clock_i _00689_ \atbs_core_0.sc_noc_generator_0.counter_value[3]\ _13989_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[4]$_DFFE_PP0P_  clock_i _00690_ \atbs_core_0.sc_noc_generator_0.counter_value[4]\ _13988_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[5]$_DFFE_PP0P_  clock_i _00691_ \atbs_core_0.sc_noc_generator_0.counter_value[5]\ _13987_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[6]$_DFFE_PP0P_  clock_i _00692_ \atbs_core_0.sc_noc_generator_0.counter_value[6]\ _00034_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_0.n2160_q[7]$_DFFE_PP0P_  clock_i _00693_ \atbs_core_0.sc_noc_generator_0.counter_value[7]\ _00035_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[0]$_DFFE_PP0P_  clock_i _00694_ \atbs_core_0.sc_noc_generator_1.counter_value[0]\ _13986_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[1]$_DFFE_PP0P_  clock_i _00695_ \atbs_core_0.sc_noc_generator_1.counter_value[1]\ _13985_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[2]$_DFFE_PP0P_  clock_i _00696_ \atbs_core_0.sc_noc_generator_1.counter_value[2]\ _13984_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[3]$_DFFE_PP0P_  clock_i _00697_ \atbs_core_0.sc_noc_generator_1.counter_value[3]\ _13983_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[4]$_DFFE_PP0P_  clock_i _00698_ \atbs_core_0.sc_noc_generator_1.counter_value[4]\ _13982_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[5]$_DFFE_PP0P_  clock_i _00699_ \atbs_core_0.sc_noc_generator_1.counter_value[5]\ _13981_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[6]$_DFFE_PP0P_  clock_i _00700_ \atbs_core_0.sc_noc_generator_1.counter_value[6]\ _00032_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_1.n2160_q[7]$_DFFE_PP0P_  clock_i _00701_ \atbs_core_0.sc_noc_generator_1.counter_value[7]\ _00033_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[0]$_DFFE_PP0P_  clock_i _00702_ \atbs_core_0.sc_noc_generator_2.counter_value[0]\ _13980_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[1]$_DFFE_PP0P_  clock_i _00703_ \atbs_core_0.sc_noc_generator_2.counter_value[1]\ _13979_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[2]$_DFFE_PP0P_  clock_i _00704_ \atbs_core_0.sc_noc_generator_2.counter_value[2]\ _13978_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[3]$_DFFE_PP0P_  clock_i _00705_ \atbs_core_0.sc_noc_generator_2.counter_value[3]\ _13977_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[4]$_DFFE_PP0P_  clock_i _00706_ \atbs_core_0.sc_noc_generator_2.counter_value[4]\ _13976_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[5]$_DFFE_PP0P_  clock_i _00707_ \atbs_core_0.sc_noc_generator_2.counter_value[5]\ _13975_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[6]$_DFFE_PP0P_  clock_i _00708_ \atbs_core_0.sc_noc_generator_2.counter_value[6]\ _00030_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_2.n2160_q[7]$_DFFE_PP0P_  clock_i _00709_ \atbs_core_0.sc_noc_generator_2.counter_value[7]\ _00031_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[0]$_DFFE_PP0P_  clock_i _00710_ \atbs_core_0.sc_noc_generator_3.counter_value[0]\ _13974_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[10]$_DFFE_PP0P_  clock_i _00711_ \atbs_core_0.sc_noc_generator_3.counter_value[10]\ _00029_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[1]$_DFFE_PP0P_  clock_i _00712_ \atbs_core_0.sc_noc_generator_3.counter_value[1]\ _13973_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[2]$_DFFE_PP0P_  clock_i _00713_ \atbs_core_0.sc_noc_generator_3.counter_value[2]\ _13972_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[3]$_DFFE_PP0P_  clock_i _00714_ \atbs_core_0.sc_noc_generator_3.counter_value[3]\ _13971_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[4]$_DFFE_PP0P_  clock_i _00715_ \atbs_core_0.sc_noc_generator_3.counter_value[4]\ _13970_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[5]$_DFFE_PP0P_  clock_i _00716_ \atbs_core_0.sc_noc_generator_3.counter_value[5]\ _13969_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[6]$_DFFE_PP0P_  clock_i _00717_ \atbs_core_0.sc_noc_generator_3.counter_value[6]\ _13968_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[7]$_DFFE_PP0P_  clock_i _00718_ \atbs_core_0.sc_noc_generator_3.counter_value[7]\ _13967_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[8]$_DFFE_PP0P_  clock_i _00719_ \atbs_core_0.sc_noc_generator_3.counter_value[8]\ _13966_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sc_noc_generator_3.n2200_q[9]$_DFFE_PP0P_  clock_i _00720_ \atbs_core_0.sc_noc_generator_3.counter_value[9]\ _00028_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1593_q$_DFF_PP0_  clock_i spike_o \atbs_core_0.spike_detector_0.hold_spike\ _00053_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1594_q$_DFFE_PP0P_  clock_i _00721_ \atbs_core_0.spike_detector_0.lock_detection\ _13965_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1595_q$_DFFE_PP0P_  clock_i _00722_ \atbs_core_0.spike_detector_0.n1595_q\ _13964_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1596_q$_DFFE_PP0P_  clock_i _00723_ \atbs_core_0.spike_detector_0.lower_is_changing\ _13963_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_detector_0.n1597_q$_DFF_PP0_  clock_i \atbs_core_0.spike_detector_0.n1583_o\ \atbs_core_0.spike_detector_0.is_changing\ _13962_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[0]$_DFFE_PP0P_  clock_i _00724_ \atbs_core_0.encoded_spike[0]\ _13961_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[10]$_DFFE_PP0P_  clock_i _00725_ \atbs_core_0.encoded_spike[10]\ _13960_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[11]$_DFFE_PP0P_  clock_i _00726_ \atbs_core_0.encoded_spike[11]\ _13959_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[12]$_DFFE_PP0P_  clock_i _00727_ \atbs_core_0.encoded_spike[12]\ _13958_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[13]$_DFFE_PP0P_  clock_i _00728_ \atbs_core_0.encoded_spike[13]\ _13957_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[14]$_DFFE_PP0P_  clock_i _00729_ \atbs_core_0.encoded_spike[14]\ _13956_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[15]$_DFFE_PP0P_  clock_i _00730_ \atbs_core_0.encoded_spike[15]\ _13955_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[16]$_DFFE_PP0P_  clock_i _00731_ \atbs_core_0.encoded_spike[16]\ _13954_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[17]$_DFFE_PP0P_  clock_i _00732_ \atbs_core_0.encoded_spike[17]\ _13953_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[18]$_DFFE_PP0P_  clock_i _00733_ \atbs_core_0.encoded_spike[18]\ _13952_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[1]$_DFFE_PP0P_  clock_i _00734_ \atbs_core_0.encoded_spike[1]\ _13951_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[2]$_DFFE_PP0P_  clock_i _00735_ \atbs_core_0.encoded_spike[2]\ _13950_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[3]$_DFFE_PP0P_  clock_i _00736_ \atbs_core_0.encoded_spike[3]\ _13949_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[4]$_DFFE_PP0P_  clock_i _00737_ \atbs_core_0.encoded_spike[4]\ _13948_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[5]$_DFFE_PP0P_  clock_i _00738_ \atbs_core_0.encoded_spike[5]\ _13947_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[6]$_DFFE_PP0P_  clock_i _00739_ \atbs_core_0.encoded_spike[6]\ _13946_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[7]$_DFFE_PP0P_  clock_i _00740_ \atbs_core_0.encoded_spike[7]\ _13945_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[8]$_DFFE_PP0P_  clock_i _00741_ \atbs_core_0.encoded_spike[8]\ _13944_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2270_q[9]$_DFFE_PP0P_  clock_i _00742_ \atbs_core_0.encoded_spike[9]\ _13943_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2271_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n2265_o\ \atbs_core_0.encoded_spike_strb\ _13942_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2272_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n2244_o\ \atbs_core_0.spike_encoder_0.delayed_spike_strb\ _13941_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_encoder_0.n2273_q$_DFF_PP0_  clock_i \atbs_core_0.spike_encoder_0.n2250_o\ \atbs_core_0.spike_encoder_0.delayed_spike\ _13940_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[0]$_DFFE_PP0P_  clock_i _00743_ \atbs_core_0.spike_memory_0.n2358_o[0]\ _13939_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1000]$_DFFE_PP0P_  clock_i _00744_ \atbs_core_0.spike_memory_0.n2410_o[12]\ _13938_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1001]$_DFFE_PP0P_  clock_i _00745_ \atbs_core_0.spike_memory_0.n2410_o[13]\ _13937_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1002]$_DFFE_PP0P_  clock_i _00746_ \atbs_core_0.spike_memory_0.n2410_o[14]\ _13936_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1003]$_DFFE_PP0P_  clock_i _00747_ \atbs_core_0.spike_memory_0.n2410_o[15]\ _13935_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1004]$_DFFE_PP0P_  clock_i _00748_ \atbs_core_0.spike_memory_0.n2410_o[16]\ _13934_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1005]$_DFFE_PP0P_  clock_i _00749_ \atbs_core_0.spike_memory_0.n2410_o[17]\ _13933_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1006]$_DFFE_PP0P_  clock_i _00750_ \atbs_core_0.spike_memory_0.n2410_o[18]\ _13932_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1007]$_DFFE_PP0P_  clock_i _00751_ \atbs_core_0.spike_memory_0.n2411_o[0]\ _13931_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1008]$_DFFE_PP0P_  clock_i _00752_ \atbs_core_0.spike_memory_0.n2411_o[1]\ _13930_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1009]$_DFFE_PP0P_  clock_i _00753_ \atbs_core_0.spike_memory_0.n2411_o[2]\ _13929_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[100]$_DFFE_PP0P_  clock_i _00754_ \atbs_core_0.spike_memory_0.n2363_o[5]\ _13928_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1010]$_DFFE_PP0P_  clock_i _00755_ \atbs_core_0.spike_memory_0.n2411_o[3]\ _13927_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1011]$_DFFE_PP0P_  clock_i _00756_ \atbs_core_0.spike_memory_0.n2411_o[4]\ _13926_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1012]$_DFFE_PP0P_  clock_i _00757_ \atbs_core_0.spike_memory_0.n2411_o[5]\ _13925_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1013]$_DFFE_PP0P_  clock_i _00758_ \atbs_core_0.spike_memory_0.n2411_o[6]\ _13924_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1014]$_DFFE_PP0P_  clock_i _00759_ \atbs_core_0.spike_memory_0.n2411_o[7]\ _13923_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1015]$_DFFE_PP0P_  clock_i _00760_ \atbs_core_0.spike_memory_0.n2411_o[8]\ _13922_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1016]$_DFFE_PP0P_  clock_i _00761_ \atbs_core_0.spike_memory_0.n2411_o[9]\ _13921_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1017]$_DFFE_PP0P_  clock_i _00762_ \atbs_core_0.spike_memory_0.n2411_o[10]\ _13920_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1018]$_DFFE_PP0P_  clock_i _00763_ \atbs_core_0.spike_memory_0.n2411_o[11]\ _13919_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1019]$_DFFE_PP0P_  clock_i _00764_ \atbs_core_0.spike_memory_0.n2411_o[12]\ _13918_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[101]$_DFFE_PP0P_  clock_i _00765_ \atbs_core_0.spike_memory_0.n2363_o[6]\ _13917_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1020]$_DFFE_PP0P_  clock_i _00766_ \atbs_core_0.spike_memory_0.n2411_o[13]\ _13916_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1021]$_DFFE_PP0P_  clock_i _00767_ \atbs_core_0.spike_memory_0.n2411_o[14]\ _13915_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1022]$_DFFE_PP0P_  clock_i _00768_ \atbs_core_0.spike_memory_0.n2411_o[15]\ _13914_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1023]$_DFFE_PP0P_  clock_i _00769_ \atbs_core_0.spike_memory_0.n2411_o[16]\ _13913_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1024]$_DFFE_PP0P_  clock_i _00770_ \atbs_core_0.spike_memory_0.n2411_o[17]\ _13912_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1025]$_DFFE_PP0P_  clock_i _00771_ \atbs_core_0.spike_memory_0.n2411_o[18]\ _13911_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1026]$_DFFE_PP0P_  clock_i _00772_ \atbs_core_0.spike_memory_0.n2412_o[0]\ _13910_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1027]$_DFFE_PP0P_  clock_i _00773_ \atbs_core_0.spike_memory_0.n2412_o[1]\ _13909_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1028]$_DFFE_PP0P_  clock_i _00774_ \atbs_core_0.spike_memory_0.n2412_o[2]\ _13908_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1029]$_DFFE_PP0P_  clock_i _00775_ \atbs_core_0.spike_memory_0.n2412_o[3]\ _13907_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[102]$_DFFE_PP0P_  clock_i _00776_ \atbs_core_0.spike_memory_0.n2363_o[7]\ _13906_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1030]$_DFFE_PP0P_  clock_i _00777_ \atbs_core_0.spike_memory_0.n2412_o[4]\ _13905_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1031]$_DFFE_PP0P_  clock_i _00778_ \atbs_core_0.spike_memory_0.n2412_o[5]\ _13904_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1032]$_DFFE_PP0P_  clock_i _00779_ \atbs_core_0.spike_memory_0.n2412_o[6]\ _13903_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1033]$_DFFE_PP0P_  clock_i _00780_ \atbs_core_0.spike_memory_0.n2412_o[7]\ _13902_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1034]$_DFFE_PP0P_  clock_i _00781_ \atbs_core_0.spike_memory_0.n2412_o[8]\ _13901_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1035]$_DFFE_PP0P_  clock_i _00782_ \atbs_core_0.spike_memory_0.n2412_o[9]\ _13900_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1036]$_DFFE_PP0P_  clock_i _00783_ \atbs_core_0.spike_memory_0.n2412_o[10]\ _13899_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1037]$_DFFE_PP0P_  clock_i _00784_ \atbs_core_0.spike_memory_0.n2412_o[11]\ _13898_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1038]$_DFFE_PP0P_  clock_i _00785_ \atbs_core_0.spike_memory_0.n2412_o[12]\ _13897_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1039]$_DFFE_PP0P_  clock_i _00786_ \atbs_core_0.spike_memory_0.n2412_o[13]\ _13896_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[103]$_DFFE_PP0P_  clock_i _00787_ \atbs_core_0.spike_memory_0.n2363_o[8]\ _13895_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1040]$_DFFE_PP0P_  clock_i _00788_ \atbs_core_0.spike_memory_0.n2412_o[14]\ _13894_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1041]$_DFFE_PP0P_  clock_i _00789_ \atbs_core_0.spike_memory_0.n2412_o[15]\ _13893_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1042]$_DFFE_PP0P_  clock_i _00790_ \atbs_core_0.spike_memory_0.n2412_o[16]\ _13892_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1043]$_DFFE_PP0P_  clock_i _00791_ \atbs_core_0.spike_memory_0.n2412_o[17]\ _13891_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1044]$_DFFE_PP0P_  clock_i _00792_ \atbs_core_0.spike_memory_0.n2412_o[18]\ _13890_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1045]$_DFFE_PP0P_  clock_i _00793_ \atbs_core_0.spike_memory_0.n2413_o[0]\ _13889_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1046]$_DFFE_PP0P_  clock_i _00794_ \atbs_core_0.spike_memory_0.n2413_o[1]\ _13888_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1047]$_DFFE_PP0P_  clock_i _00795_ \atbs_core_0.spike_memory_0.n2413_o[2]\ _13887_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1048]$_DFFE_PP0P_  clock_i _00796_ \atbs_core_0.spike_memory_0.n2413_o[3]\ _13886_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1049]$_DFFE_PP0P_  clock_i _00797_ \atbs_core_0.spike_memory_0.n2413_o[4]\ _13885_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[104]$_DFFE_PP0P_  clock_i _00798_ \atbs_core_0.spike_memory_0.n2363_o[9]\ _13884_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1050]$_DFFE_PP0P_  clock_i _00799_ \atbs_core_0.spike_memory_0.n2413_o[5]\ _13883_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1051]$_DFFE_PP0P_  clock_i _00800_ \atbs_core_0.spike_memory_0.n2413_o[6]\ _13882_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1052]$_DFFE_PP0P_  clock_i _00801_ \atbs_core_0.spike_memory_0.n2413_o[7]\ _13881_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1053]$_DFFE_PP0P_  clock_i _00802_ \atbs_core_0.spike_memory_0.n2413_o[8]\ _13880_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1054]$_DFFE_PP0P_  clock_i _00803_ \atbs_core_0.spike_memory_0.n2413_o[9]\ _13879_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1055]$_DFFE_PP0P_  clock_i _00804_ \atbs_core_0.spike_memory_0.n2413_o[10]\ _13878_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1056]$_DFFE_PP0P_  clock_i _00805_ \atbs_core_0.spike_memory_0.n2413_o[11]\ _13877_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1057]$_DFFE_PP0P_  clock_i _00806_ \atbs_core_0.spike_memory_0.n2413_o[12]\ _13876_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1058]$_DFFE_PP0P_  clock_i _00807_ \atbs_core_0.spike_memory_0.n2413_o[13]\ _13875_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1059]$_DFFE_PP0P_  clock_i _00808_ \atbs_core_0.spike_memory_0.n2413_o[14]\ _13874_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[105]$_DFFE_PP0P_  clock_i _00809_ \atbs_core_0.spike_memory_0.n2363_o[10]\ _13873_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1060]$_DFFE_PP0P_  clock_i _00810_ \atbs_core_0.spike_memory_0.n2413_o[15]\ _13872_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1061]$_DFFE_PP0P_  clock_i _00811_ \atbs_core_0.spike_memory_0.n2413_o[16]\ _13871_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1062]$_DFFE_PP0P_  clock_i _00812_ \atbs_core_0.spike_memory_0.n2413_o[17]\ _13870_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1063]$_DFFE_PP0P_  clock_i _00813_ \atbs_core_0.spike_memory_0.n2413_o[18]\ _13869_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1064]$_DFFE_PP0P_  clock_i _00814_ \atbs_core_0.spike_memory_0.n2414_o[0]\ _13868_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1065]$_DFFE_PP0P_  clock_i _00815_ \atbs_core_0.spike_memory_0.n2414_o[1]\ _13867_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1066]$_DFFE_PP0P_  clock_i _00816_ \atbs_core_0.spike_memory_0.n2414_o[2]\ _13866_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1067]$_DFFE_PP0P_  clock_i _00817_ \atbs_core_0.spike_memory_0.n2414_o[3]\ _13865_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1068]$_DFFE_PP0P_  clock_i _00818_ \atbs_core_0.spike_memory_0.n2414_o[4]\ _13864_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1069]$_DFFE_PP0P_  clock_i _00819_ \atbs_core_0.spike_memory_0.n2414_o[5]\ _13863_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[106]$_DFFE_PP0P_  clock_i _00820_ \atbs_core_0.spike_memory_0.n2363_o[11]\ _13862_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1070]$_DFFE_PP0P_  clock_i _00821_ \atbs_core_0.spike_memory_0.n2414_o[6]\ _13861_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1071]$_DFFE_PP0P_  clock_i _00822_ \atbs_core_0.spike_memory_0.n2414_o[7]\ _13860_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1072]$_DFFE_PP0P_  clock_i _00823_ \atbs_core_0.spike_memory_0.n2414_o[8]\ _13859_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1073]$_DFFE_PP0P_  clock_i _00824_ \atbs_core_0.spike_memory_0.n2414_o[9]\ _13858_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1074]$_DFFE_PP0P_  clock_i _00825_ \atbs_core_0.spike_memory_0.n2414_o[10]\ _13857_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1075]$_DFFE_PP0P_  clock_i _00826_ \atbs_core_0.spike_memory_0.n2414_o[11]\ _13856_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1076]$_DFFE_PP0P_  clock_i _00827_ \atbs_core_0.spike_memory_0.n2414_o[12]\ _13855_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1077]$_DFFE_PP0P_  clock_i _00828_ \atbs_core_0.spike_memory_0.n2414_o[13]\ _13854_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1078]$_DFFE_PP0P_  clock_i _00829_ \atbs_core_0.spike_memory_0.n2414_o[14]\ _13853_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1079]$_DFFE_PP0P_  clock_i _00830_ \atbs_core_0.spike_memory_0.n2414_o[15]\ _13852_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[107]$_DFFE_PP0P_  clock_i _00831_ \atbs_core_0.spike_memory_0.n2363_o[12]\ _13851_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1080]$_DFFE_PP0P_  clock_i _00832_ \atbs_core_0.spike_memory_0.n2414_o[16]\ _13850_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1081]$_DFFE_PP0P_  clock_i _00833_ \atbs_core_0.spike_memory_0.n2414_o[17]\ _13849_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1082]$_DFFE_PP0P_  clock_i _00834_ \atbs_core_0.spike_memory_0.n2414_o[18]\ _13848_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1083]$_DFFE_PP0P_  clock_i _00835_ \atbs_core_0.spike_memory_0.n2415_o[0]\ _13847_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1084]$_DFFE_PP0P_  clock_i _00836_ \atbs_core_0.spike_memory_0.n2415_o[1]\ _13846_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1085]$_DFFE_PP0P_  clock_i _00837_ \atbs_core_0.spike_memory_0.n2415_o[2]\ _13845_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1086]$_DFFE_PP0P_  clock_i _00838_ \atbs_core_0.spike_memory_0.n2415_o[3]\ _13844_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1087]$_DFFE_PP0P_  clock_i _00839_ \atbs_core_0.spike_memory_0.n2415_o[4]\ _13843_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1088]$_DFFE_PP0P_  clock_i _00840_ \atbs_core_0.spike_memory_0.n2415_o[5]\ _13842_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1089]$_DFFE_PP0P_  clock_i _00841_ \atbs_core_0.spike_memory_0.n2415_o[6]\ _13841_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[108]$_DFFE_PP0P_  clock_i _00842_ \atbs_core_0.spike_memory_0.n2363_o[13]\ _13840_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1090]$_DFFE_PP0P_  clock_i _00843_ \atbs_core_0.spike_memory_0.n2415_o[7]\ _13839_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1091]$_DFFE_PP0P_  clock_i _00844_ \atbs_core_0.spike_memory_0.n2415_o[8]\ _13838_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1092]$_DFFE_PP0P_  clock_i _00845_ \atbs_core_0.spike_memory_0.n2415_o[9]\ _13837_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1093]$_DFFE_PP0P_  clock_i _00846_ \atbs_core_0.spike_memory_0.n2415_o[10]\ _13836_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1094]$_DFFE_PP0P_  clock_i _00847_ \atbs_core_0.spike_memory_0.n2415_o[11]\ _13835_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1095]$_DFFE_PP0P_  clock_i _00848_ \atbs_core_0.spike_memory_0.n2415_o[12]\ _13834_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1096]$_DFFE_PP0P_  clock_i _00849_ \atbs_core_0.spike_memory_0.n2415_o[13]\ _13833_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1097]$_DFFE_PP0P_  clock_i _00850_ \atbs_core_0.spike_memory_0.n2415_o[14]\ _13832_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1098]$_DFFE_PP0P_  clock_i _00851_ \atbs_core_0.spike_memory_0.n2415_o[15]\ _13831_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1099]$_DFFE_PP0P_  clock_i _00852_ \atbs_core_0.spike_memory_0.n2415_o[16]\ _13830_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[109]$_DFFE_PP0P_  clock_i _00853_ \atbs_core_0.spike_memory_0.n2363_o[14]\ _13829_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[10]$_DFFE_PP0P_  clock_i _00854_ \atbs_core_0.spike_memory_0.n2358_o[10]\ _13828_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1100]$_DFFE_PP0P_  clock_i _00855_ \atbs_core_0.spike_memory_0.n2415_o[17]\ _13827_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1101]$_DFFE_PP0P_  clock_i _00856_ \atbs_core_0.spike_memory_0.n2415_o[18]\ _13826_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1102]$_DFFE_PP0P_  clock_i _00857_ \atbs_core_0.spike_memory_0.n2416_o[0]\ _13825_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1103]$_DFFE_PP0P_  clock_i _00858_ \atbs_core_0.spike_memory_0.n2416_o[1]\ _13824_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1104]$_DFFE_PP0P_  clock_i _00859_ \atbs_core_0.spike_memory_0.n2416_o[2]\ _13823_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1105]$_DFFE_PP0P_  clock_i _00860_ \atbs_core_0.spike_memory_0.n2416_o[3]\ _13822_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1106]$_DFFE_PP0P_  clock_i _00861_ \atbs_core_0.spike_memory_0.n2416_o[4]\ _13821_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1107]$_DFFE_PP0P_  clock_i _00862_ \atbs_core_0.spike_memory_0.n2416_o[5]\ _13820_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1108]$_DFFE_PP0P_  clock_i _00863_ \atbs_core_0.spike_memory_0.n2416_o[6]\ _13819_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1109]$_DFFE_PP0P_  clock_i _00864_ \atbs_core_0.spike_memory_0.n2416_o[7]\ _13818_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[110]$_DFFE_PP0P_  clock_i _00865_ \atbs_core_0.spike_memory_0.n2363_o[15]\ _13817_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1110]$_DFFE_PP0P_  clock_i _00866_ \atbs_core_0.spike_memory_0.n2416_o[8]\ _13816_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1111]$_DFFE_PP0P_  clock_i _00867_ \atbs_core_0.spike_memory_0.n2416_o[9]\ _13815_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1112]$_DFFE_PP0P_  clock_i _00868_ \atbs_core_0.spike_memory_0.n2416_o[10]\ _13814_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1113]$_DFFE_PP0P_  clock_i _00869_ \atbs_core_0.spike_memory_0.n2416_o[11]\ _13813_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1114]$_DFFE_PP0P_  clock_i _00870_ \atbs_core_0.spike_memory_0.n2416_o[12]\ _13812_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1115]$_DFFE_PP0P_  clock_i _00871_ \atbs_core_0.spike_memory_0.n2416_o[13]\ _13811_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1116]$_DFFE_PP0P_  clock_i _00872_ \atbs_core_0.spike_memory_0.n2416_o[14]\ _13810_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1117]$_DFFE_PP0P_  clock_i _00873_ \atbs_core_0.spike_memory_0.n2416_o[15]\ _13809_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1118]$_DFFE_PP0P_  clock_i _00874_ \atbs_core_0.spike_memory_0.n2416_o[16]\ _13808_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1119]$_DFFE_PP0P_  clock_i _00875_ \atbs_core_0.spike_memory_0.n2416_o[17]\ _13807_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[111]$_DFFE_PP0P_  clock_i _00876_ \atbs_core_0.spike_memory_0.n2363_o[16]\ _13806_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1120]$_DFFE_PP0P_  clock_i _00877_ \atbs_core_0.spike_memory_0.n2416_o[18]\ _13805_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1121]$_DFFE_PP0P_  clock_i _00878_ \atbs_core_0.spike_memory_0.n2417_o[0]\ _13804_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1122]$_DFFE_PP0P_  clock_i _00879_ \atbs_core_0.spike_memory_0.n2417_o[1]\ _13803_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1123]$_DFFE_PP0P_  clock_i _00880_ \atbs_core_0.spike_memory_0.n2417_o[2]\ _13802_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1124]$_DFFE_PP0P_  clock_i _00881_ \atbs_core_0.spike_memory_0.n2417_o[3]\ _13801_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1125]$_DFFE_PP0P_  clock_i _00882_ \atbs_core_0.spike_memory_0.n2417_o[4]\ _13800_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1126]$_DFFE_PP0P_  clock_i _00883_ \atbs_core_0.spike_memory_0.n2417_o[5]\ _13799_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1127]$_DFFE_PP0P_  clock_i _00884_ \atbs_core_0.spike_memory_0.n2417_o[6]\ _13798_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1128]$_DFFE_PP0P_  clock_i _00885_ \atbs_core_0.spike_memory_0.n2417_o[7]\ _13797_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1129]$_DFFE_PP0P_  clock_i _00886_ \atbs_core_0.spike_memory_0.n2417_o[8]\ _13796_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[112]$_DFFE_PP0P_  clock_i _00887_ \atbs_core_0.spike_memory_0.n2363_o[17]\ _13795_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1130]$_DFFE_PP0P_  clock_i _00888_ \atbs_core_0.spike_memory_0.n2417_o[9]\ _13794_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1131]$_DFFE_PP0P_  clock_i _00889_ \atbs_core_0.spike_memory_0.n2417_o[10]\ _13793_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1132]$_DFFE_PP0P_  clock_i _00890_ \atbs_core_0.spike_memory_0.n2417_o[11]\ _13792_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1133]$_DFFE_PP0P_  clock_i _00891_ \atbs_core_0.spike_memory_0.n2417_o[12]\ _13791_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1134]$_DFFE_PP0P_  clock_i _00892_ \atbs_core_0.spike_memory_0.n2417_o[13]\ _13790_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1135]$_DFFE_PP0P_  clock_i _00893_ \atbs_core_0.spike_memory_0.n2417_o[14]\ _13789_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1136]$_DFFE_PP0P_  clock_i _00894_ \atbs_core_0.spike_memory_0.n2417_o[15]\ _13788_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1137]$_DFFE_PP0P_  clock_i _00895_ \atbs_core_0.spike_memory_0.n2417_o[16]\ _13787_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1138]$_DFFE_PP0P_  clock_i _00896_ \atbs_core_0.spike_memory_0.n2417_o[17]\ _13786_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1139]$_DFFE_PP0P_  clock_i _00897_ \atbs_core_0.spike_memory_0.n2417_o[18]\ _13785_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[113]$_DFFE_PP0P_  clock_i _00898_ \atbs_core_0.spike_memory_0.n2363_o[18]\ _13784_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1140]$_DFFE_PP0P_  clock_i _00899_ \atbs_core_0.spike_memory_0.n2418_o[0]\ _13783_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1141]$_DFFE_PP0P_  clock_i _00900_ \atbs_core_0.spike_memory_0.n2418_o[1]\ _13782_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1142]$_DFFE_PP0P_  clock_i _00901_ \atbs_core_0.spike_memory_0.n2418_o[2]\ _13781_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1143]$_DFFE_PP0P_  clock_i _00902_ \atbs_core_0.spike_memory_0.n2418_o[3]\ _13780_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1144]$_DFFE_PP0P_  clock_i _00903_ \atbs_core_0.spike_memory_0.n2418_o[4]\ _13779_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1145]$_DFFE_PP0P_  clock_i _00904_ \atbs_core_0.spike_memory_0.n2418_o[5]\ _13778_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1146]$_DFFE_PP0P_  clock_i _00905_ \atbs_core_0.spike_memory_0.n2418_o[6]\ _13777_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1147]$_DFFE_PP0P_  clock_i _00906_ \atbs_core_0.spike_memory_0.n2418_o[7]\ _13776_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1148]$_DFFE_PP0P_  clock_i _00907_ \atbs_core_0.spike_memory_0.n2418_o[8]\ _13775_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1149]$_DFFE_PP0P_  clock_i _00908_ \atbs_core_0.spike_memory_0.n2418_o[9]\ _13774_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[114]$_DFFE_PP0P_  clock_i _00909_ \atbs_core_0.spike_memory_0.n2364_o[0]\ _13773_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1150]$_DFFE_PP0P_  clock_i _00910_ \atbs_core_0.spike_memory_0.n2418_o[10]\ _13772_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1151]$_DFFE_PP0P_  clock_i _00911_ \atbs_core_0.spike_memory_0.n2418_o[11]\ _13771_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1152]$_DFFE_PP0P_  clock_i _00912_ \atbs_core_0.spike_memory_0.n2418_o[12]\ _13770_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1153]$_DFFE_PP0P_  clock_i _00913_ \atbs_core_0.spike_memory_0.n2418_o[13]\ _13769_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1154]$_DFFE_PP0P_  clock_i _00914_ \atbs_core_0.spike_memory_0.n2418_o[14]\ _13768_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1155]$_DFFE_PP0P_  clock_i _00915_ \atbs_core_0.spike_memory_0.n2418_o[15]\ _13767_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1156]$_DFFE_PP0P_  clock_i _00916_ \atbs_core_0.spike_memory_0.n2418_o[16]\ _13766_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1157]$_DFFE_PP0P_  clock_i _00917_ \atbs_core_0.spike_memory_0.n2418_o[17]\ _13765_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1158]$_DFFE_PP0P_  clock_i _00918_ \atbs_core_0.spike_memory_0.n2418_o[18]\ _13764_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1159]$_DFFE_PP0P_  clock_i _00919_ \atbs_core_0.spike_memory_0.n2419_o[0]\ _13763_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[115]$_DFFE_PP0P_  clock_i _00920_ \atbs_core_0.spike_memory_0.n2364_o[1]\ _13762_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1160]$_DFFE_PP0P_  clock_i _00921_ \atbs_core_0.spike_memory_0.n2419_o[1]\ _13761_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1161]$_DFFE_PP0P_  clock_i _00922_ \atbs_core_0.spike_memory_0.n2419_o[2]\ _13760_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1162]$_DFFE_PP0P_  clock_i _00923_ \atbs_core_0.spike_memory_0.n2419_o[3]\ _13759_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1163]$_DFFE_PP0P_  clock_i _00924_ \atbs_core_0.spike_memory_0.n2419_o[4]\ _13758_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1164]$_DFFE_PP0P_  clock_i _00925_ \atbs_core_0.spike_memory_0.n2419_o[5]\ _13757_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1165]$_DFFE_PP0P_  clock_i _00926_ \atbs_core_0.spike_memory_0.n2419_o[6]\ _13756_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1166]$_DFFE_PP0P_  clock_i _00927_ \atbs_core_0.spike_memory_0.n2419_o[7]\ _13755_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1167]$_DFFE_PP0P_  clock_i _00928_ \atbs_core_0.spike_memory_0.n2419_o[8]\ _13754_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1168]$_DFFE_PP0P_  clock_i _00929_ \atbs_core_0.spike_memory_0.n2419_o[9]\ _13753_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1169]$_DFFE_PP0P_  clock_i _00930_ \atbs_core_0.spike_memory_0.n2419_o[10]\ _13752_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[116]$_DFFE_PP0P_  clock_i _00931_ \atbs_core_0.spike_memory_0.n2364_o[2]\ _13751_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1170]$_DFFE_PP0P_  clock_i _00932_ \atbs_core_0.spike_memory_0.n2419_o[11]\ _13750_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1171]$_DFFE_PP0P_  clock_i _00933_ \atbs_core_0.spike_memory_0.n2419_o[12]\ _13749_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1172]$_DFFE_PP0P_  clock_i _00934_ \atbs_core_0.spike_memory_0.n2419_o[13]\ _13748_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1173]$_DFFE_PP0P_  clock_i _00935_ \atbs_core_0.spike_memory_0.n2419_o[14]\ _13747_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1174]$_DFFE_PP0P_  clock_i _00936_ \atbs_core_0.spike_memory_0.n2419_o[15]\ _13746_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1175]$_DFFE_PP0P_  clock_i _00937_ \atbs_core_0.spike_memory_0.n2419_o[16]\ _13745_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1176]$_DFFE_PP0P_  clock_i _00938_ \atbs_core_0.spike_memory_0.n2419_o[17]\ _13744_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1177]$_DFFE_PP0P_  clock_i _00939_ \atbs_core_0.spike_memory_0.n2419_o[18]\ _13743_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1178]$_DFFE_PP0P_  clock_i _00940_ \atbs_core_0.spike_memory_0.n2420_o[0]\ _13742_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1179]$_DFFE_PP0P_  clock_i _00941_ \atbs_core_0.spike_memory_0.n2420_o[1]\ _13741_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[117]$_DFFE_PP0P_  clock_i _00942_ \atbs_core_0.spike_memory_0.n2364_o[3]\ _13740_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1180]$_DFFE_PP0P_  clock_i _00943_ \atbs_core_0.spike_memory_0.n2420_o[2]\ _13739_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1181]$_DFFE_PP0P_  clock_i _00944_ \atbs_core_0.spike_memory_0.n2420_o[3]\ _13738_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1182]$_DFFE_PP0P_  clock_i _00945_ \atbs_core_0.spike_memory_0.n2420_o[4]\ _13737_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1183]$_DFFE_PP0P_  clock_i _00946_ \atbs_core_0.spike_memory_0.n2420_o[5]\ _13736_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1184]$_DFFE_PP0P_  clock_i _00947_ \atbs_core_0.spike_memory_0.n2420_o[6]\ _13735_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1185]$_DFFE_PP0P_  clock_i _00948_ \atbs_core_0.spike_memory_0.n2420_o[7]\ _13734_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1186]$_DFFE_PP0P_  clock_i _00949_ \atbs_core_0.spike_memory_0.n2420_o[8]\ _13733_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1187]$_DFFE_PP0P_  clock_i _00950_ \atbs_core_0.spike_memory_0.n2420_o[9]\ _13732_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1188]$_DFFE_PP0P_  clock_i _00951_ \atbs_core_0.spike_memory_0.n2420_o[10]\ _13731_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1189]$_DFFE_PP0P_  clock_i _00952_ \atbs_core_0.spike_memory_0.n2420_o[11]\ _13730_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[118]$_DFFE_PP0P_  clock_i _00953_ \atbs_core_0.spike_memory_0.n2364_o[4]\ _13729_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1190]$_DFFE_PP0P_  clock_i _00954_ \atbs_core_0.spike_memory_0.n2420_o[12]\ _13728_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1191]$_DFFE_PP0P_  clock_i _00955_ \atbs_core_0.spike_memory_0.n2420_o[13]\ _13727_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1192]$_DFFE_PP0P_  clock_i _00956_ \atbs_core_0.spike_memory_0.n2420_o[14]\ _13726_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1193]$_DFFE_PP0P_  clock_i _00957_ \atbs_core_0.spike_memory_0.n2420_o[15]\ _13725_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1194]$_DFFE_PP0P_  clock_i _00958_ \atbs_core_0.spike_memory_0.n2420_o[16]\ _13724_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1195]$_DFFE_PP0P_  clock_i _00959_ \atbs_core_0.spike_memory_0.n2420_o[17]\ _13723_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1196]$_DFFE_PP0P_  clock_i _00960_ \atbs_core_0.spike_memory_0.n2420_o[18]\ _13722_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1197]$_DFFE_PP0P_  clock_i _00961_ \atbs_core_0.spike_memory_0.n2436_q[1197]\ _13721_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1198]$_DFFE_PP0P_  clock_i _00962_ \atbs_core_0.spike_memory_0.n2436_q[1198]\ _13720_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1199]$_DFFE_PP0P_  clock_i _00963_ \atbs_core_0.spike_memory_0.n2436_q[1199]\ _13719_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[119]$_DFFE_PP0P_  clock_i _00964_ \atbs_core_0.spike_memory_0.n2364_o[5]\ _13718_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[11]$_DFFE_PP0P_  clock_i _00965_ \atbs_core_0.spike_memory_0.n2358_o[11]\ _13717_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1200]$_DFFE_PP0P_  clock_i _00966_ \atbs_core_0.spike_memory_0.n2436_q[1200]\ _13716_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1201]$_DFFE_PP0P_  clock_i _00967_ \atbs_core_0.spike_memory_0.n2436_q[1201]\ _13715_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1202]$_DFFE_PP0P_  clock_i _00968_ \atbs_core_0.spike_memory_0.n2436_q[1202]\ _13714_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1203]$_DFFE_PP0P_  clock_i _00969_ \atbs_core_0.spike_memory_0.n2436_q[1203]\ _13713_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1204]$_DFFE_PP0P_  clock_i _00970_ \atbs_core_0.spike_memory_0.n2436_q[1204]\ _13712_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1205]$_DFFE_PP0P_  clock_i _00971_ \atbs_core_0.spike_memory_0.n2436_q[1205]\ _13711_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1206]$_DFFE_PP0P_  clock_i _00972_ \atbs_core_0.spike_memory_0.n2436_q[1206]\ _13710_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1207]$_DFFE_PP0P_  clock_i _00973_ \atbs_core_0.spike_memory_0.n2436_q[1207]\ _13709_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1208]$_DFFE_PP0P_  clock_i _00974_ \atbs_core_0.spike_memory_0.n2436_q[1208]\ _13708_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1209]$_DFFE_PP0P_  clock_i _00975_ \atbs_core_0.spike_memory_0.n2436_q[1209]\ _13707_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[120]$_DFFE_PP0P_  clock_i _00976_ \atbs_core_0.spike_memory_0.n2364_o[6]\ _13706_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1210]$_DFFE_PP0P_  clock_i _00977_ \atbs_core_0.spike_memory_0.n2436_q[1210]\ _13705_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1211]$_DFFE_PP0P_  clock_i _00978_ \atbs_core_0.spike_memory_0.n2436_q[1211]\ _13704_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1212]$_DFFE_PP0P_  clock_i _00979_ \atbs_core_0.spike_memory_0.n2436_q[1212]\ _13703_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1213]$_DFFE_PP0P_  clock_i _00980_ \atbs_core_0.spike_memory_0.n2436_q[1213]\ _13702_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1214]$_DFFE_PP0P_  clock_i _00981_ \atbs_core_0.spike_memory_0.n2436_q[1214]\ _13701_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1215]$_DFFE_PP0P_  clock_i _00982_ \atbs_core_0.spike_memory_0.n2436_q[1215]\ _13700_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[121]$_DFFE_PP0P_  clock_i _00983_ \atbs_core_0.spike_memory_0.n2364_o[7]\ _13699_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[122]$_DFFE_PP0P_  clock_i _00984_ \atbs_core_0.spike_memory_0.n2364_o[8]\ _13698_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[123]$_DFFE_PP0P_  clock_i _00985_ \atbs_core_0.spike_memory_0.n2364_o[9]\ _13697_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[124]$_DFFE_PP0P_  clock_i _00986_ \atbs_core_0.spike_memory_0.n2364_o[10]\ _13696_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[125]$_DFFE_PP0P_  clock_i _00987_ \atbs_core_0.spike_memory_0.n2364_o[11]\ _13695_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[126]$_DFFE_PP0P_  clock_i _00988_ \atbs_core_0.spike_memory_0.n2364_o[12]\ _13694_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[127]$_DFFE_PP0P_  clock_i _00989_ \atbs_core_0.spike_memory_0.n2364_o[13]\ _13693_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[128]$_DFFE_PP0P_  clock_i _00990_ \atbs_core_0.spike_memory_0.n2364_o[14]\ _13692_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[129]$_DFFE_PP0P_  clock_i _00991_ \atbs_core_0.spike_memory_0.n2364_o[15]\ _13691_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[12]$_DFFE_PP0P_  clock_i _00992_ \atbs_core_0.spike_memory_0.n2358_o[12]\ _13690_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[130]$_DFFE_PP0P_  clock_i _00993_ \atbs_core_0.spike_memory_0.n2364_o[16]\ _13689_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[131]$_DFFE_PP0P_  clock_i _00994_ \atbs_core_0.spike_memory_0.n2364_o[17]\ _13688_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[132]$_DFFE_PP0P_  clock_i _00995_ \atbs_core_0.spike_memory_0.n2364_o[18]\ _13687_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[133]$_DFFE_PP0P_  clock_i _00996_ \atbs_core_0.spike_memory_0.n2365_o[0]\ _13686_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[134]$_DFFE_PP0P_  clock_i _00997_ \atbs_core_0.spike_memory_0.n2365_o[1]\ _13685_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[135]$_DFFE_PP0P_  clock_i _00998_ \atbs_core_0.spike_memory_0.n2365_o[2]\ _13684_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[136]$_DFFE_PP0P_  clock_i _00999_ \atbs_core_0.spike_memory_0.n2365_o[3]\ _13683_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[137]$_DFFE_PP0P_  clock_i _01000_ \atbs_core_0.spike_memory_0.n2365_o[4]\ _13682_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[138]$_DFFE_PP0P_  clock_i _01001_ \atbs_core_0.spike_memory_0.n2365_o[5]\ _13681_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[139]$_DFFE_PP0P_  clock_i _01002_ \atbs_core_0.spike_memory_0.n2365_o[6]\ _13680_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[13]$_DFFE_PP0P_  clock_i _01003_ \atbs_core_0.spike_memory_0.n2358_o[13]\ _13679_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[140]$_DFFE_PP0P_  clock_i _01004_ \atbs_core_0.spike_memory_0.n2365_o[7]\ _13678_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[141]$_DFFE_PP0P_  clock_i _01005_ \atbs_core_0.spike_memory_0.n2365_o[8]\ _13677_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[142]$_DFFE_PP0P_  clock_i _01006_ \atbs_core_0.spike_memory_0.n2365_o[9]\ _13676_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[143]$_DFFE_PP0P_  clock_i _01007_ \atbs_core_0.spike_memory_0.n2365_o[10]\ _13675_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[144]$_DFFE_PP0P_  clock_i _01008_ \atbs_core_0.spike_memory_0.n2365_o[11]\ _13674_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[145]$_DFFE_PP0P_  clock_i _01009_ \atbs_core_0.spike_memory_0.n2365_o[12]\ _13673_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[146]$_DFFE_PP0P_  clock_i _01010_ \atbs_core_0.spike_memory_0.n2365_o[13]\ _13672_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[147]$_DFFE_PP0P_  clock_i _01011_ \atbs_core_0.spike_memory_0.n2365_o[14]\ _13671_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[148]$_DFFE_PP0P_  clock_i _01012_ \atbs_core_0.spike_memory_0.n2365_o[15]\ _13670_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[149]$_DFFE_PP0P_  clock_i _01013_ \atbs_core_0.spike_memory_0.n2365_o[16]\ _13669_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[14]$_DFFE_PP0P_  clock_i _01014_ \atbs_core_0.spike_memory_0.n2358_o[14]\ _13668_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[150]$_DFFE_PP0P_  clock_i _01015_ \atbs_core_0.spike_memory_0.n2365_o[17]\ _13667_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[151]$_DFFE_PP0P_  clock_i _01016_ \atbs_core_0.spike_memory_0.n2365_o[18]\ _13666_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[152]$_DFFE_PP0P_  clock_i _01017_ \atbs_core_0.spike_memory_0.n2366_o[0]\ _13665_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[153]$_DFFE_PP0P_  clock_i _01018_ \atbs_core_0.spike_memory_0.n2366_o[1]\ _13664_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[154]$_DFFE_PP0P_  clock_i _01019_ \atbs_core_0.spike_memory_0.n2366_o[2]\ _13663_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[155]$_DFFE_PP0P_  clock_i _01020_ \atbs_core_0.spike_memory_0.n2366_o[3]\ _13662_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[156]$_DFFE_PP0P_  clock_i _01021_ \atbs_core_0.spike_memory_0.n2366_o[4]\ _13661_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[157]$_DFFE_PP0P_  clock_i _01022_ \atbs_core_0.spike_memory_0.n2366_o[5]\ _13660_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[158]$_DFFE_PP0P_  clock_i _01023_ \atbs_core_0.spike_memory_0.n2366_o[6]\ _13659_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[159]$_DFFE_PP0P_  clock_i _01024_ \atbs_core_0.spike_memory_0.n2366_o[7]\ _13658_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[15]$_DFFE_PP0P_  clock_i _01025_ \atbs_core_0.spike_memory_0.n2358_o[15]\ _13657_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[160]$_DFFE_PP0P_  clock_i _01026_ \atbs_core_0.spike_memory_0.n2366_o[8]\ _13656_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[161]$_DFFE_PP0P_  clock_i _01027_ \atbs_core_0.spike_memory_0.n2366_o[9]\ _13655_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[162]$_DFFE_PP0P_  clock_i _01028_ \atbs_core_0.spike_memory_0.n2366_o[10]\ _13654_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[163]$_DFFE_PP0P_  clock_i _01029_ \atbs_core_0.spike_memory_0.n2366_o[11]\ _13653_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[164]$_DFFE_PP0P_  clock_i _01030_ \atbs_core_0.spike_memory_0.n2366_o[12]\ _13652_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[165]$_DFFE_PP0P_  clock_i _01031_ \atbs_core_0.spike_memory_0.n2366_o[13]\ _13651_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[166]$_DFFE_PP0P_  clock_i _01032_ \atbs_core_0.spike_memory_0.n2366_o[14]\ _13650_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[167]$_DFFE_PP0P_  clock_i _01033_ \atbs_core_0.spike_memory_0.n2366_o[15]\ _13649_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[168]$_DFFE_PP0P_  clock_i _01034_ \atbs_core_0.spike_memory_0.n2366_o[16]\ _13648_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[169]$_DFFE_PP0P_  clock_i _01035_ \atbs_core_0.spike_memory_0.n2366_o[17]\ _13647_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[16]$_DFFE_PP0P_  clock_i _01036_ \atbs_core_0.spike_memory_0.n2358_o[16]\ _13646_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[170]$_DFFE_PP0P_  clock_i _01037_ \atbs_core_0.spike_memory_0.n2366_o[18]\ _13645_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[171]$_DFFE_PP0P_  clock_i _01038_ \atbs_core_0.spike_memory_0.n2367_o[0]\ _13644_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[172]$_DFFE_PP0P_  clock_i _01039_ \atbs_core_0.spike_memory_0.n2367_o[1]\ _13643_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[173]$_DFFE_PP0P_  clock_i _01040_ \atbs_core_0.spike_memory_0.n2367_o[2]\ _13642_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[174]$_DFFE_PP0P_  clock_i _01041_ \atbs_core_0.spike_memory_0.n2367_o[3]\ _13641_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[175]$_DFFE_PP0P_  clock_i _01042_ \atbs_core_0.spike_memory_0.n2367_o[4]\ _13640_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[176]$_DFFE_PP0P_  clock_i _01043_ \atbs_core_0.spike_memory_0.n2367_o[5]\ _13639_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[177]$_DFFE_PP0P_  clock_i _01044_ \atbs_core_0.spike_memory_0.n2367_o[6]\ _13638_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[178]$_DFFE_PP0P_  clock_i _01045_ \atbs_core_0.spike_memory_0.n2367_o[7]\ _13637_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[179]$_DFFE_PP0P_  clock_i _01046_ \atbs_core_0.spike_memory_0.n2367_o[8]\ _13636_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[17]$_DFFE_PP0P_  clock_i _01047_ \atbs_core_0.spike_memory_0.n2358_o[17]\ _13635_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[180]$_DFFE_PP0P_  clock_i _01048_ \atbs_core_0.spike_memory_0.n2367_o[9]\ _13634_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[181]$_DFFE_PP0P_  clock_i _01049_ \atbs_core_0.spike_memory_0.n2367_o[10]\ _13633_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[182]$_DFFE_PP0P_  clock_i _01050_ \atbs_core_0.spike_memory_0.n2367_o[11]\ _13632_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[183]$_DFFE_PP0P_  clock_i _01051_ \atbs_core_0.spike_memory_0.n2367_o[12]\ _13631_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[184]$_DFFE_PP0P_  clock_i _01052_ \atbs_core_0.spike_memory_0.n2367_o[13]\ _13630_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[185]$_DFFE_PP0P_  clock_i _01053_ \atbs_core_0.spike_memory_0.n2367_o[14]\ _13629_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[186]$_DFFE_PP0P_  clock_i _01054_ \atbs_core_0.spike_memory_0.n2367_o[15]\ _13628_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[187]$_DFFE_PP0P_  clock_i _01055_ \atbs_core_0.spike_memory_0.n2367_o[16]\ _13627_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[188]$_DFFE_PP0P_  clock_i _01056_ \atbs_core_0.spike_memory_0.n2367_o[17]\ _13626_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[189]$_DFFE_PP0P_  clock_i _01057_ \atbs_core_0.spike_memory_0.n2367_o[18]\ _13625_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[18]$_DFFE_PP0P_  clock_i _01058_ \atbs_core_0.spike_memory_0.n2358_o[18]\ _13624_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[190]$_DFFE_PP0P_  clock_i _01059_ \atbs_core_0.spike_memory_0.n2368_o[0]\ _13623_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[191]$_DFFE_PP0P_  clock_i _01060_ \atbs_core_0.spike_memory_0.n2368_o[1]\ _13622_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[192]$_DFFE_PP0P_  clock_i _01061_ \atbs_core_0.spike_memory_0.n2368_o[2]\ _13621_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[193]$_DFFE_PP0P_  clock_i _01062_ \atbs_core_0.spike_memory_0.n2368_o[3]\ _13620_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[194]$_DFFE_PP0P_  clock_i _01063_ \atbs_core_0.spike_memory_0.n2368_o[4]\ _13619_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[195]$_DFFE_PP0P_  clock_i _01064_ \atbs_core_0.spike_memory_0.n2368_o[5]\ _13618_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[196]$_DFFE_PP0P_  clock_i _01065_ \atbs_core_0.spike_memory_0.n2368_o[6]\ _13617_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[197]$_DFFE_PP0P_  clock_i _01066_ \atbs_core_0.spike_memory_0.n2368_o[7]\ _13616_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[198]$_DFFE_PP0P_  clock_i _01067_ \atbs_core_0.spike_memory_0.n2368_o[8]\ _13615_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[199]$_DFFE_PP0P_  clock_i _01068_ \atbs_core_0.spike_memory_0.n2368_o[9]\ _13614_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[19]$_DFFE_PP0P_  clock_i _01069_ \atbs_core_0.spike_memory_0.n2359_o[0]\ _13613_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[1]$_DFFE_PP0P_  clock_i _01070_ \atbs_core_0.spike_memory_0.n2358_o[1]\ _13612_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[200]$_DFFE_PP0P_  clock_i _01071_ \atbs_core_0.spike_memory_0.n2368_o[10]\ _13611_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[201]$_DFFE_PP0P_  clock_i _01072_ \atbs_core_0.spike_memory_0.n2368_o[11]\ _13610_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[202]$_DFFE_PP0P_  clock_i _01073_ \atbs_core_0.spike_memory_0.n2368_o[12]\ _13609_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[203]$_DFFE_PP0P_  clock_i _01074_ \atbs_core_0.spike_memory_0.n2368_o[13]\ _13608_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[204]$_DFFE_PP0P_  clock_i _01075_ \atbs_core_0.spike_memory_0.n2368_o[14]\ _13607_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[205]$_DFFE_PP0P_  clock_i _01076_ \atbs_core_0.spike_memory_0.n2368_o[15]\ _13606_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[206]$_DFFE_PP0P_  clock_i _01077_ \atbs_core_0.spike_memory_0.n2368_o[16]\ _13605_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[207]$_DFFE_PP0P_  clock_i _01078_ \atbs_core_0.spike_memory_0.n2368_o[17]\ _13604_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[208]$_DFFE_PP0P_  clock_i _01079_ \atbs_core_0.spike_memory_0.n2368_o[18]\ _13603_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[209]$_DFFE_PP0P_  clock_i _01080_ \atbs_core_0.spike_memory_0.n2369_o[0]\ _13602_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[20]$_DFFE_PP0P_  clock_i _01081_ \atbs_core_0.spike_memory_0.n2359_o[1]\ _13601_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[210]$_DFFE_PP0P_  clock_i _01082_ \atbs_core_0.spike_memory_0.n2369_o[1]\ _13600_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[211]$_DFFE_PP0P_  clock_i _01083_ \atbs_core_0.spike_memory_0.n2369_o[2]\ _13599_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[212]$_DFFE_PP0P_  clock_i _01084_ \atbs_core_0.spike_memory_0.n2369_o[3]\ _13598_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[213]$_DFFE_PP0P_  clock_i _01085_ \atbs_core_0.spike_memory_0.n2369_o[4]\ _13597_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[214]$_DFFE_PP0P_  clock_i _01086_ \atbs_core_0.spike_memory_0.n2369_o[5]\ _13596_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[215]$_DFFE_PP0P_  clock_i _01087_ \atbs_core_0.spike_memory_0.n2369_o[6]\ _13595_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[216]$_DFFE_PP0P_  clock_i _01088_ \atbs_core_0.spike_memory_0.n2369_o[7]\ _13594_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[217]$_DFFE_PP0P_  clock_i _01089_ \atbs_core_0.spike_memory_0.n2369_o[8]\ _13593_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[218]$_DFFE_PP0P_  clock_i _01090_ \atbs_core_0.spike_memory_0.n2369_o[9]\ _13592_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[219]$_DFFE_PP0P_  clock_i _01091_ \atbs_core_0.spike_memory_0.n2369_o[10]\ _13591_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[21]$_DFFE_PP0P_  clock_i _01092_ \atbs_core_0.spike_memory_0.n2359_o[2]\ _13590_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[220]$_DFFE_PP0P_  clock_i _01093_ \atbs_core_0.spike_memory_0.n2369_o[11]\ _13589_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[221]$_DFFE_PP0P_  clock_i _01094_ \atbs_core_0.spike_memory_0.n2369_o[12]\ _13588_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[222]$_DFFE_PP0P_  clock_i _01095_ \atbs_core_0.spike_memory_0.n2369_o[13]\ _13587_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[223]$_DFFE_PP0P_  clock_i _01096_ \atbs_core_0.spike_memory_0.n2369_o[14]\ _13586_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[224]$_DFFE_PP0P_  clock_i _01097_ \atbs_core_0.spike_memory_0.n2369_o[15]\ _13585_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[225]$_DFFE_PP0P_  clock_i _01098_ \atbs_core_0.spike_memory_0.n2369_o[16]\ _13584_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[226]$_DFFE_PP0P_  clock_i _01099_ \atbs_core_0.spike_memory_0.n2369_o[17]\ _13583_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[227]$_DFFE_PP0P_  clock_i _01100_ \atbs_core_0.spike_memory_0.n2369_o[18]\ _13582_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[228]$_DFFE_PP0P_  clock_i _01101_ \atbs_core_0.spike_memory_0.n2370_o[0]\ _13581_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[229]$_DFFE_PP0P_  clock_i _01102_ \atbs_core_0.spike_memory_0.n2370_o[1]\ _13580_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[22]$_DFFE_PP0P_  clock_i _01103_ \atbs_core_0.spike_memory_0.n2359_o[3]\ _13579_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[230]$_DFFE_PP0P_  clock_i _01104_ \atbs_core_0.spike_memory_0.n2370_o[2]\ _13578_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[231]$_DFFE_PP0P_  clock_i _01105_ \atbs_core_0.spike_memory_0.n2370_o[3]\ _13577_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[232]$_DFFE_PP0P_  clock_i _01106_ \atbs_core_0.spike_memory_0.n2370_o[4]\ _13576_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[233]$_DFFE_PP0P_  clock_i _01107_ \atbs_core_0.spike_memory_0.n2370_o[5]\ _13575_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[234]$_DFFE_PP0P_  clock_i _01108_ \atbs_core_0.spike_memory_0.n2370_o[6]\ _13574_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[235]$_DFFE_PP0P_  clock_i _01109_ \atbs_core_0.spike_memory_0.n2370_o[7]\ _13573_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[236]$_DFFE_PP0P_  clock_i _01110_ \atbs_core_0.spike_memory_0.n2370_o[8]\ _13572_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[237]$_DFFE_PP0P_  clock_i _01111_ \atbs_core_0.spike_memory_0.n2370_o[9]\ _13571_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[238]$_DFFE_PP0P_  clock_i _01112_ \atbs_core_0.spike_memory_0.n2370_o[10]\ _13570_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[239]$_DFFE_PP0P_  clock_i _01113_ \atbs_core_0.spike_memory_0.n2370_o[11]\ _13569_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[23]$_DFFE_PP0P_  clock_i _01114_ \atbs_core_0.spike_memory_0.n2359_o[4]\ _13568_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[240]$_DFFE_PP0P_  clock_i _01115_ \atbs_core_0.spike_memory_0.n2370_o[12]\ _13567_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[241]$_DFFE_PP0P_  clock_i _01116_ \atbs_core_0.spike_memory_0.n2370_o[13]\ _13566_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[242]$_DFFE_PP0P_  clock_i _01117_ \atbs_core_0.spike_memory_0.n2370_o[14]\ _13565_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[243]$_DFFE_PP0P_  clock_i _01118_ \atbs_core_0.spike_memory_0.n2370_o[15]\ _13564_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[244]$_DFFE_PP0P_  clock_i _01119_ \atbs_core_0.spike_memory_0.n2370_o[16]\ _13563_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[245]$_DFFE_PP0P_  clock_i _01120_ \atbs_core_0.spike_memory_0.n2370_o[17]\ _13562_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[246]$_DFFE_PP0P_  clock_i _01121_ \atbs_core_0.spike_memory_0.n2370_o[18]\ _13561_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[247]$_DFFE_PP0P_  clock_i _01122_ \atbs_core_0.spike_memory_0.n2371_o[0]\ _13560_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[248]$_DFFE_PP0P_  clock_i _01123_ \atbs_core_0.spike_memory_0.n2371_o[1]\ _13559_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[249]$_DFFE_PP0P_  clock_i _01124_ \atbs_core_0.spike_memory_0.n2371_o[2]\ _13558_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[24]$_DFFE_PP0P_  clock_i _01125_ \atbs_core_0.spike_memory_0.n2359_o[5]\ _13557_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[250]$_DFFE_PP0P_  clock_i _01126_ \atbs_core_0.spike_memory_0.n2371_o[3]\ _13556_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[251]$_DFFE_PP0P_  clock_i _01127_ \atbs_core_0.spike_memory_0.n2371_o[4]\ _13555_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[252]$_DFFE_PP0P_  clock_i _01128_ \atbs_core_0.spike_memory_0.n2371_o[5]\ _13554_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[253]$_DFFE_PP0P_  clock_i _01129_ \atbs_core_0.spike_memory_0.n2371_o[6]\ _13553_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[254]$_DFFE_PP0P_  clock_i _01130_ \atbs_core_0.spike_memory_0.n2371_o[7]\ _13552_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[255]$_DFFE_PP0P_  clock_i _01131_ \atbs_core_0.spike_memory_0.n2371_o[8]\ _13551_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[256]$_DFFE_PP0P_  clock_i _01132_ \atbs_core_0.spike_memory_0.n2371_o[9]\ _13550_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[257]$_DFFE_PP0P_  clock_i _01133_ \atbs_core_0.spike_memory_0.n2371_o[10]\ _13549_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[258]$_DFFE_PP0P_  clock_i _01134_ \atbs_core_0.spike_memory_0.n2371_o[11]\ _13548_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[259]$_DFFE_PP0P_  clock_i _01135_ \atbs_core_0.spike_memory_0.n2371_o[12]\ _13547_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[25]$_DFFE_PP0P_  clock_i _01136_ \atbs_core_0.spike_memory_0.n2359_o[6]\ _13546_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[260]$_DFFE_PP0P_  clock_i _01137_ \atbs_core_0.spike_memory_0.n2371_o[13]\ _13545_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[261]$_DFFE_PP0P_  clock_i _01138_ \atbs_core_0.spike_memory_0.n2371_o[14]\ _13544_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[262]$_DFFE_PP0P_  clock_i _01139_ \atbs_core_0.spike_memory_0.n2371_o[15]\ _13543_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[263]$_DFFE_PP0P_  clock_i _01140_ \atbs_core_0.spike_memory_0.n2371_o[16]\ _13542_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[264]$_DFFE_PP0P_  clock_i _01141_ \atbs_core_0.spike_memory_0.n2371_o[17]\ _13541_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[265]$_DFFE_PP0P_  clock_i _01142_ \atbs_core_0.spike_memory_0.n2371_o[18]\ _13540_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[266]$_DFFE_PP0P_  clock_i _01143_ \atbs_core_0.spike_memory_0.n2372_o[0]\ _13539_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[267]$_DFFE_PP0P_  clock_i _01144_ \atbs_core_0.spike_memory_0.n2372_o[1]\ _13538_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[268]$_DFFE_PP0P_  clock_i _01145_ \atbs_core_0.spike_memory_0.n2372_o[2]\ _13537_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[269]$_DFFE_PP0P_  clock_i _01146_ \atbs_core_0.spike_memory_0.n2372_o[3]\ _13536_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[26]$_DFFE_PP0P_  clock_i _01147_ \atbs_core_0.spike_memory_0.n2359_o[7]\ _13535_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[270]$_DFFE_PP0P_  clock_i _01148_ \atbs_core_0.spike_memory_0.n2372_o[4]\ _13534_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[271]$_DFFE_PP0P_  clock_i _01149_ \atbs_core_0.spike_memory_0.n2372_o[5]\ _13533_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[272]$_DFFE_PP0P_  clock_i _01150_ \atbs_core_0.spike_memory_0.n2372_o[6]\ _13532_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[273]$_DFFE_PP0P_  clock_i _01151_ \atbs_core_0.spike_memory_0.n2372_o[7]\ _13531_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[274]$_DFFE_PP0P_  clock_i _01152_ \atbs_core_0.spike_memory_0.n2372_o[8]\ _13530_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[275]$_DFFE_PP0P_  clock_i _01153_ \atbs_core_0.spike_memory_0.n2372_o[9]\ _13529_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[276]$_DFFE_PP0P_  clock_i _01154_ \atbs_core_0.spike_memory_0.n2372_o[10]\ _13528_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[277]$_DFFE_PP0P_  clock_i _01155_ \atbs_core_0.spike_memory_0.n2372_o[11]\ _13527_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[278]$_DFFE_PP0P_  clock_i _01156_ \atbs_core_0.spike_memory_0.n2372_o[12]\ _13526_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[279]$_DFFE_PP0P_  clock_i _01157_ \atbs_core_0.spike_memory_0.n2372_o[13]\ _13525_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[27]$_DFFE_PP0P_  clock_i _01158_ \atbs_core_0.spike_memory_0.n2359_o[8]\ _13524_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[280]$_DFFE_PP0P_  clock_i _01159_ \atbs_core_0.spike_memory_0.n2372_o[14]\ _13523_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[281]$_DFFE_PP0P_  clock_i _01160_ \atbs_core_0.spike_memory_0.n2372_o[15]\ _13522_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[282]$_DFFE_PP0P_  clock_i _01161_ \atbs_core_0.spike_memory_0.n2372_o[16]\ _13521_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[283]$_DFFE_PP0P_  clock_i _01162_ \atbs_core_0.spike_memory_0.n2372_o[17]\ _13520_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[284]$_DFFE_PP0P_  clock_i _01163_ \atbs_core_0.spike_memory_0.n2372_o[18]\ _13519_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[285]$_DFFE_PP0P_  clock_i _01164_ \atbs_core_0.spike_memory_0.n2373_o[0]\ _13518_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[286]$_DFFE_PP0P_  clock_i _01165_ \atbs_core_0.spike_memory_0.n2373_o[1]\ _13517_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[287]$_DFFE_PP0P_  clock_i _01166_ \atbs_core_0.spike_memory_0.n2373_o[2]\ _13516_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[288]$_DFFE_PP0P_  clock_i _01167_ \atbs_core_0.spike_memory_0.n2373_o[3]\ _13515_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[289]$_DFFE_PP0P_  clock_i _01168_ \atbs_core_0.spike_memory_0.n2373_o[4]\ _13514_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[28]$_DFFE_PP0P_  clock_i _01169_ \atbs_core_0.spike_memory_0.n2359_o[9]\ _13513_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[290]$_DFFE_PP0P_  clock_i _01170_ \atbs_core_0.spike_memory_0.n2373_o[5]\ _13512_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[291]$_DFFE_PP0P_  clock_i _01171_ \atbs_core_0.spike_memory_0.n2373_o[6]\ _13511_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[292]$_DFFE_PP0P_  clock_i _01172_ \atbs_core_0.spike_memory_0.n2373_o[7]\ _13510_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[293]$_DFFE_PP0P_  clock_i _01173_ \atbs_core_0.spike_memory_0.n2373_o[8]\ _13509_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[294]$_DFFE_PP0P_  clock_i _01174_ \atbs_core_0.spike_memory_0.n2373_o[9]\ _13508_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[295]$_DFFE_PP0P_  clock_i _01175_ \atbs_core_0.spike_memory_0.n2373_o[10]\ _13507_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[296]$_DFFE_PP0P_  clock_i _01176_ \atbs_core_0.spike_memory_0.n2373_o[11]\ _13506_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[297]$_DFFE_PP0P_  clock_i _01177_ \atbs_core_0.spike_memory_0.n2373_o[12]\ _13505_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[298]$_DFFE_PP0P_  clock_i _01178_ \atbs_core_0.spike_memory_0.n2373_o[13]\ _13504_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[299]$_DFFE_PP0P_  clock_i _01179_ \atbs_core_0.spike_memory_0.n2373_o[14]\ _13503_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[29]$_DFFE_PP0P_  clock_i _01180_ \atbs_core_0.spike_memory_0.n2359_o[10]\ _13502_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[2]$_DFFE_PP0P_  clock_i _01181_ \atbs_core_0.spike_memory_0.n2358_o[2]\ _13501_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[300]$_DFFE_PP0P_  clock_i _01182_ \atbs_core_0.spike_memory_0.n2373_o[15]\ _13500_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[301]$_DFFE_PP0P_  clock_i _01183_ \atbs_core_0.spike_memory_0.n2373_o[16]\ _13499_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[302]$_DFFE_PP0P_  clock_i _01184_ \atbs_core_0.spike_memory_0.n2373_o[17]\ _13498_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[303]$_DFFE_PP0P_  clock_i _01185_ \atbs_core_0.spike_memory_0.n2373_o[18]\ _13497_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[304]$_DFFE_PP0P_  clock_i _01186_ \atbs_core_0.spike_memory_0.n2374_o[0]\ _00112_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[305]$_DFFE_PP0P_  clock_i _01187_ \atbs_core_0.spike_memory_0.n2374_o[1]\ _00115_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[306]$_DFFE_PP0P_  clock_i _01188_ \atbs_core_0.spike_memory_0.n2374_o[2]\ _00118_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[307]$_DFFE_PP0P_  clock_i _01189_ \atbs_core_0.spike_memory_0.n2374_o[3]\ _00121_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[308]$_DFFE_PP0P_  clock_i _01190_ \atbs_core_0.spike_memory_0.n2374_o[4]\ _00124_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[309]$_DFFE_PP0P_  clock_i _01191_ \atbs_core_0.spike_memory_0.n2374_o[5]\ _00127_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[30]$_DFFE_PP0P_  clock_i _01192_ \atbs_core_0.spike_memory_0.n2359_o[11]\ _13496_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[310]$_DFFE_PP0P_  clock_i _01193_ \atbs_core_0.spike_memory_0.n2374_o[6]\ _00130_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[311]$_DFFE_PP0P_  clock_i _01194_ \atbs_core_0.spike_memory_0.n2374_o[7]\ _00133_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[312]$_DFFE_PP0P_  clock_i _01195_ \atbs_core_0.spike_memory_0.n2374_o[8]\ _00136_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[313]$_DFFE_PP0P_  clock_i _01196_ \atbs_core_0.spike_memory_0.n2374_o[9]\ _00139_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[314]$_DFFE_PP0P_  clock_i _01197_ \atbs_core_0.spike_memory_0.n2374_o[10]\ _00142_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[315]$_DFFE_PP0P_  clock_i _01198_ \atbs_core_0.spike_memory_0.n2374_o[11]\ _00145_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[316]$_DFFE_PP0P_  clock_i _01199_ \atbs_core_0.spike_memory_0.n2374_o[12]\ _00148_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[317]$_DFFE_PP0P_  clock_i _01200_ \atbs_core_0.spike_memory_0.n2374_o[13]\ _00006_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[318]$_DFFE_PP0P_  clock_i _01201_ \atbs_core_0.spike_memory_0.n2374_o[14]\ _00009_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[319]$_DFFE_PP0P_  clock_i _01202_ \atbs_core_0.spike_memory_0.n2374_o[15]\ _00012_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[31]$_DFFE_PP0P_  clock_i _01203_ \atbs_core_0.spike_memory_0.n2359_o[12]\ _13495_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[320]$_DFFE_PP0P_  clock_i _01204_ \atbs_core_0.spike_memory_0.n2374_o[16]\ _00015_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[321]$_DFFE_PP0P_  clock_i _01205_ \atbs_core_0.spike_memory_0.n2374_o[17]\ _00018_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[322]$_DFFE_PP0P_  clock_i _01206_ \atbs_core_0.spike_memory_0.n2374_o[18]\ _00021_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[323]$_DFFE_PP0P_  clock_i _01207_ \atbs_core_0.spike_memory_0.n2375_o[0]\ _13494_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[324]$_DFFE_PP0P_  clock_i _01208_ \atbs_core_0.spike_memory_0.n2375_o[1]\ _13493_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[325]$_DFFE_PP0P_  clock_i _01209_ \atbs_core_0.spike_memory_0.n2375_o[2]\ _13492_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[326]$_DFFE_PP0P_  clock_i _01210_ \atbs_core_0.spike_memory_0.n2375_o[3]\ _13491_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[327]$_DFFE_PP0P_  clock_i _01211_ \atbs_core_0.spike_memory_0.n2375_o[4]\ _13490_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[328]$_DFFE_PP0P_  clock_i _01212_ \atbs_core_0.spike_memory_0.n2375_o[5]\ _13489_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[329]$_DFFE_PP0P_  clock_i _01213_ \atbs_core_0.spike_memory_0.n2375_o[6]\ _13488_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[32]$_DFFE_PP0P_  clock_i _01214_ \atbs_core_0.spike_memory_0.n2359_o[13]\ _13487_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[330]$_DFFE_PP0P_  clock_i _01215_ \atbs_core_0.spike_memory_0.n2375_o[7]\ _13486_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[331]$_DFFE_PP0P_  clock_i _01216_ \atbs_core_0.spike_memory_0.n2375_o[8]\ _13485_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[332]$_DFFE_PP0P_  clock_i _01217_ \atbs_core_0.spike_memory_0.n2375_o[9]\ _13484_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[333]$_DFFE_PP0P_  clock_i _01218_ \atbs_core_0.spike_memory_0.n2375_o[10]\ _13483_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[334]$_DFFE_PP0P_  clock_i _01219_ \atbs_core_0.spike_memory_0.n2375_o[11]\ _13482_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[335]$_DFFE_PP0P_  clock_i _01220_ \atbs_core_0.spike_memory_0.n2375_o[12]\ _13481_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[336]$_DFFE_PP0P_  clock_i _01221_ \atbs_core_0.spike_memory_0.n2375_o[13]\ _13480_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[337]$_DFFE_PP0P_  clock_i _01222_ \atbs_core_0.spike_memory_0.n2375_o[14]\ _13479_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[338]$_DFFE_PP0P_  clock_i _01223_ \atbs_core_0.spike_memory_0.n2375_o[15]\ _13478_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[339]$_DFFE_PP0P_  clock_i _01224_ \atbs_core_0.spike_memory_0.n2375_o[16]\ _13477_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[33]$_DFFE_PP0P_  clock_i _01225_ \atbs_core_0.spike_memory_0.n2359_o[14]\ _13476_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[340]$_DFFE_PP0P_  clock_i _01226_ \atbs_core_0.spike_memory_0.n2375_o[17]\ _13475_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[341]$_DFFE_PP0P_  clock_i _01227_ \atbs_core_0.spike_memory_0.n2375_o[18]\ _13474_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[342]$_DFFE_PP0P_  clock_i _01228_ \atbs_core_0.spike_memory_0.n2376_o[0]\ _13473_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[343]$_DFFE_PP0P_  clock_i _01229_ \atbs_core_0.spike_memory_0.n2376_o[1]\ _13472_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[344]$_DFFE_PP0P_  clock_i _01230_ \atbs_core_0.spike_memory_0.n2376_o[2]\ _13471_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[345]$_DFFE_PP0P_  clock_i _01231_ \atbs_core_0.spike_memory_0.n2376_o[3]\ _13470_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[346]$_DFFE_PP0P_  clock_i _01232_ \atbs_core_0.spike_memory_0.n2376_o[4]\ _13469_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[347]$_DFFE_PP0P_  clock_i _01233_ \atbs_core_0.spike_memory_0.n2376_o[5]\ _13468_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[348]$_DFFE_PP0P_  clock_i _01234_ \atbs_core_0.spike_memory_0.n2376_o[6]\ _13467_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[349]$_DFFE_PP0P_  clock_i _01235_ \atbs_core_0.spike_memory_0.n2376_o[7]\ _13466_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[34]$_DFFE_PP0P_  clock_i _01236_ \atbs_core_0.spike_memory_0.n2359_o[15]\ _13465_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[350]$_DFFE_PP0P_  clock_i _01237_ \atbs_core_0.spike_memory_0.n2376_o[8]\ _13464_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[351]$_DFFE_PP0P_  clock_i _01238_ \atbs_core_0.spike_memory_0.n2376_o[9]\ _13463_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[352]$_DFFE_PP0P_  clock_i _01239_ \atbs_core_0.spike_memory_0.n2376_o[10]\ _13462_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[353]$_DFFE_PP0P_  clock_i _01240_ \atbs_core_0.spike_memory_0.n2376_o[11]\ _13461_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[354]$_DFFE_PP0P_  clock_i _01241_ \atbs_core_0.spike_memory_0.n2376_o[12]\ _13460_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[355]$_DFFE_PP0P_  clock_i _01242_ \atbs_core_0.spike_memory_0.n2376_o[13]\ _13459_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[356]$_DFFE_PP0P_  clock_i _01243_ \atbs_core_0.spike_memory_0.n2376_o[14]\ _13458_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[357]$_DFFE_PP0P_  clock_i _01244_ \atbs_core_0.spike_memory_0.n2376_o[15]\ _13457_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[358]$_DFFE_PP0P_  clock_i _01245_ \atbs_core_0.spike_memory_0.n2376_o[16]\ _13456_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[359]$_DFFE_PP0P_  clock_i _01246_ \atbs_core_0.spike_memory_0.n2376_o[17]\ _13455_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[35]$_DFFE_PP0P_  clock_i _01247_ \atbs_core_0.spike_memory_0.n2359_o[16]\ _13454_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[360]$_DFFE_PP0P_  clock_i _01248_ \atbs_core_0.spike_memory_0.n2376_o[18]\ _13453_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[361]$_DFFE_PP0P_  clock_i _01249_ \atbs_core_0.spike_memory_0.n2377_o[0]\ _13452_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[362]$_DFFE_PP0P_  clock_i _01250_ \atbs_core_0.spike_memory_0.n2377_o[1]\ _13451_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[363]$_DFFE_PP0P_  clock_i _01251_ \atbs_core_0.spike_memory_0.n2377_o[2]\ _13450_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[364]$_DFFE_PP0P_  clock_i _01252_ \atbs_core_0.spike_memory_0.n2377_o[3]\ _13449_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[365]$_DFFE_PP0P_  clock_i _01253_ \atbs_core_0.spike_memory_0.n2377_o[4]\ _13448_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[366]$_DFFE_PP0P_  clock_i _01254_ \atbs_core_0.spike_memory_0.n2377_o[5]\ _13447_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[367]$_DFFE_PP0P_  clock_i _01255_ \atbs_core_0.spike_memory_0.n2377_o[6]\ _13446_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[368]$_DFFE_PP0P_  clock_i _01256_ \atbs_core_0.spike_memory_0.n2377_o[7]\ _13445_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[369]$_DFFE_PP0P_  clock_i _01257_ \atbs_core_0.spike_memory_0.n2377_o[8]\ _13444_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[36]$_DFFE_PP0P_  clock_i _01258_ \atbs_core_0.spike_memory_0.n2359_o[17]\ _13443_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[370]$_DFFE_PP0P_  clock_i _01259_ \atbs_core_0.spike_memory_0.n2377_o[9]\ _13442_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[371]$_DFFE_PP0P_  clock_i _01260_ \atbs_core_0.spike_memory_0.n2377_o[10]\ _13441_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[372]$_DFFE_PP0P_  clock_i _01261_ \atbs_core_0.spike_memory_0.n2377_o[11]\ _13440_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[373]$_DFFE_PP0P_  clock_i _01262_ \atbs_core_0.spike_memory_0.n2377_o[12]\ _13439_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[374]$_DFFE_PP0P_  clock_i _01263_ \atbs_core_0.spike_memory_0.n2377_o[13]\ _13438_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[375]$_DFFE_PP0P_  clock_i _01264_ \atbs_core_0.spike_memory_0.n2377_o[14]\ _13437_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[376]$_DFFE_PP0P_  clock_i _01265_ \atbs_core_0.spike_memory_0.n2377_o[15]\ _13436_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[377]$_DFFE_PP0P_  clock_i _01266_ \atbs_core_0.spike_memory_0.n2377_o[16]\ _13435_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[378]$_DFFE_PP0P_  clock_i _01267_ \atbs_core_0.spike_memory_0.n2377_o[17]\ _13434_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[379]$_DFFE_PP0P_  clock_i _01268_ \atbs_core_0.spike_memory_0.n2377_o[18]\ _13433_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[37]$_DFFE_PP0P_  clock_i _01269_ \atbs_core_0.spike_memory_0.n2359_o[18]\ _13432_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[380]$_DFFE_PP0P_  clock_i _01270_ \atbs_core_0.spike_memory_0.n2378_o[0]\ _13431_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[381]$_DFFE_PP0P_  clock_i _01271_ \atbs_core_0.spike_memory_0.n2378_o[1]\ _13430_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[382]$_DFFE_PP0P_  clock_i _01272_ \atbs_core_0.spike_memory_0.n2378_o[2]\ _13429_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[383]$_DFFE_PP0P_  clock_i _01273_ \atbs_core_0.spike_memory_0.n2378_o[3]\ _13428_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[384]$_DFFE_PP0P_  clock_i _01274_ \atbs_core_0.spike_memory_0.n2378_o[4]\ _13427_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[385]$_DFFE_PP0P_  clock_i _01275_ \atbs_core_0.spike_memory_0.n2378_o[5]\ _13426_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[386]$_DFFE_PP0P_  clock_i _01276_ \atbs_core_0.spike_memory_0.n2378_o[6]\ _13425_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[387]$_DFFE_PP0P_  clock_i _01277_ \atbs_core_0.spike_memory_0.n2378_o[7]\ _13424_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[388]$_DFFE_PP0P_  clock_i _01278_ \atbs_core_0.spike_memory_0.n2378_o[8]\ _13423_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[389]$_DFFE_PP0P_  clock_i _01279_ \atbs_core_0.spike_memory_0.n2378_o[9]\ _13422_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[38]$_DFFE_PP0P_  clock_i _01280_ \atbs_core_0.spike_memory_0.n2360_o[0]\ _13421_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[390]$_DFFE_PP0P_  clock_i _01281_ \atbs_core_0.spike_memory_0.n2378_o[10]\ _13420_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[391]$_DFFE_PP0P_  clock_i _01282_ \atbs_core_0.spike_memory_0.n2378_o[11]\ _13419_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[392]$_DFFE_PP0P_  clock_i _01283_ \atbs_core_0.spike_memory_0.n2378_o[12]\ _13418_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[393]$_DFFE_PP0P_  clock_i _01284_ \atbs_core_0.spike_memory_0.n2378_o[13]\ _13417_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[394]$_DFFE_PP0P_  clock_i _01285_ \atbs_core_0.spike_memory_0.n2378_o[14]\ _13416_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[395]$_DFFE_PP0P_  clock_i _01286_ \atbs_core_0.spike_memory_0.n2378_o[15]\ _13415_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[396]$_DFFE_PP0P_  clock_i _01287_ \atbs_core_0.spike_memory_0.n2378_o[16]\ _13414_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[397]$_DFFE_PP0P_  clock_i _01288_ \atbs_core_0.spike_memory_0.n2378_o[17]\ _13413_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[398]$_DFFE_PP0P_  clock_i _01289_ \atbs_core_0.spike_memory_0.n2378_o[18]\ _13412_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[399]$_DFFE_PP0P_  clock_i _01290_ \atbs_core_0.spike_memory_0.n2379_o[0]\ _13411_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[39]$_DFFE_PP0P_  clock_i _01291_ \atbs_core_0.spike_memory_0.n2360_o[1]\ _13410_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[3]$_DFFE_PP0P_  clock_i _01292_ \atbs_core_0.spike_memory_0.n2358_o[3]\ _13409_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[400]$_DFFE_PP0P_  clock_i _01293_ \atbs_core_0.spike_memory_0.n2379_o[1]\ _13408_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[401]$_DFFE_PP0P_  clock_i _01294_ \atbs_core_0.spike_memory_0.n2379_o[2]\ _13407_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[402]$_DFFE_PP0P_  clock_i _01295_ \atbs_core_0.spike_memory_0.n2379_o[3]\ _13406_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[403]$_DFFE_PP0P_  clock_i _01296_ \atbs_core_0.spike_memory_0.n2379_o[4]\ _13405_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[404]$_DFFE_PP0P_  clock_i _01297_ \atbs_core_0.spike_memory_0.n2379_o[5]\ _13404_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[405]$_DFFE_PP0P_  clock_i _01298_ \atbs_core_0.spike_memory_0.n2379_o[6]\ _13403_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[406]$_DFFE_PP0P_  clock_i _01299_ \atbs_core_0.spike_memory_0.n2379_o[7]\ _13402_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[407]$_DFFE_PP0P_  clock_i _01300_ \atbs_core_0.spike_memory_0.n2379_o[8]\ _13401_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[408]$_DFFE_PP0P_  clock_i _01301_ \atbs_core_0.spike_memory_0.n2379_o[9]\ _13400_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[409]$_DFFE_PP0P_  clock_i _01302_ \atbs_core_0.spike_memory_0.n2379_o[10]\ _13399_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[40]$_DFFE_PP0P_  clock_i _01303_ \atbs_core_0.spike_memory_0.n2360_o[2]\ _13398_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[410]$_DFFE_PP0P_  clock_i _01304_ \atbs_core_0.spike_memory_0.n2379_o[11]\ _13397_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[411]$_DFFE_PP0P_  clock_i _01305_ \atbs_core_0.spike_memory_0.n2379_o[12]\ _13396_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[412]$_DFFE_PP0P_  clock_i _01306_ \atbs_core_0.spike_memory_0.n2379_o[13]\ _13395_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[413]$_DFFE_PP0P_  clock_i _01307_ \atbs_core_0.spike_memory_0.n2379_o[14]\ _13394_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[414]$_DFFE_PP0P_  clock_i _01308_ \atbs_core_0.spike_memory_0.n2379_o[15]\ _13393_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[415]$_DFFE_PP0P_  clock_i _01309_ \atbs_core_0.spike_memory_0.n2379_o[16]\ _13392_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[416]$_DFFE_PP0P_  clock_i _01310_ \atbs_core_0.spike_memory_0.n2379_o[17]\ _13391_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[417]$_DFFE_PP0P_  clock_i _01311_ \atbs_core_0.spike_memory_0.n2379_o[18]\ _13390_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[418]$_DFFE_PP0P_  clock_i _01312_ \atbs_core_0.spike_memory_0.n2380_o[0]\ _13389_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[419]$_DFFE_PP0P_  clock_i _01313_ \atbs_core_0.spike_memory_0.n2380_o[1]\ _13388_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[41]$_DFFE_PP0P_  clock_i _01314_ \atbs_core_0.spike_memory_0.n2360_o[3]\ _13387_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[420]$_DFFE_PP0P_  clock_i _01315_ \atbs_core_0.spike_memory_0.n2380_o[2]\ _13386_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[421]$_DFFE_PP0P_  clock_i _01316_ \atbs_core_0.spike_memory_0.n2380_o[3]\ _13385_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[422]$_DFFE_PP0P_  clock_i _01317_ \atbs_core_0.spike_memory_0.n2380_o[4]\ _13384_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[423]$_DFFE_PP0P_  clock_i _01318_ \atbs_core_0.spike_memory_0.n2380_o[5]\ _13383_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[424]$_DFFE_PP0P_  clock_i _01319_ \atbs_core_0.spike_memory_0.n2380_o[6]\ _13382_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[425]$_DFFE_PP0P_  clock_i _01320_ \atbs_core_0.spike_memory_0.n2380_o[7]\ _13381_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[426]$_DFFE_PP0P_  clock_i _01321_ \atbs_core_0.spike_memory_0.n2380_o[8]\ _13380_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[427]$_DFFE_PP0P_  clock_i _01322_ \atbs_core_0.spike_memory_0.n2380_o[9]\ _13379_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[428]$_DFFE_PP0P_  clock_i _01323_ \atbs_core_0.spike_memory_0.n2380_o[10]\ _13378_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[429]$_DFFE_PP0P_  clock_i _01324_ \atbs_core_0.spike_memory_0.n2380_o[11]\ _13377_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[42]$_DFFE_PP0P_  clock_i _01325_ \atbs_core_0.spike_memory_0.n2360_o[4]\ _13376_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[430]$_DFFE_PP0P_  clock_i _01326_ \atbs_core_0.spike_memory_0.n2380_o[12]\ _13375_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[431]$_DFFE_PP0P_  clock_i _01327_ \atbs_core_0.spike_memory_0.n2380_o[13]\ _13374_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[432]$_DFFE_PP0P_  clock_i _01328_ \atbs_core_0.spike_memory_0.n2380_o[14]\ _13373_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[433]$_DFFE_PP0P_  clock_i _01329_ \atbs_core_0.spike_memory_0.n2380_o[15]\ _13372_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[434]$_DFFE_PP0P_  clock_i _01330_ \atbs_core_0.spike_memory_0.n2380_o[16]\ _13371_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[435]$_DFFE_PP0P_  clock_i _01331_ \atbs_core_0.spike_memory_0.n2380_o[17]\ _13370_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[436]$_DFFE_PP0P_  clock_i _01332_ \atbs_core_0.spike_memory_0.n2380_o[18]\ _13369_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[437]$_DFFE_PP0P_  clock_i _01333_ \atbs_core_0.spike_memory_0.n2381_o[0]\ _13368_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[438]$_DFFE_PP0P_  clock_i _01334_ \atbs_core_0.spike_memory_0.n2381_o[1]\ _13367_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[439]$_DFFE_PP0P_  clock_i _01335_ \atbs_core_0.spike_memory_0.n2381_o[2]\ _13366_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[43]$_DFFE_PP0P_  clock_i _01336_ \atbs_core_0.spike_memory_0.n2360_o[5]\ _13365_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[440]$_DFFE_PP0P_  clock_i _01337_ \atbs_core_0.spike_memory_0.n2381_o[3]\ _13364_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[441]$_DFFE_PP0P_  clock_i _01338_ \atbs_core_0.spike_memory_0.n2381_o[4]\ _13363_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[442]$_DFFE_PP0P_  clock_i _01339_ \atbs_core_0.spike_memory_0.n2381_o[5]\ _13362_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[443]$_DFFE_PP0P_  clock_i _01340_ \atbs_core_0.spike_memory_0.n2381_o[6]\ _13361_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[444]$_DFFE_PP0P_  clock_i _01341_ \atbs_core_0.spike_memory_0.n2381_o[7]\ _13360_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[445]$_DFFE_PP0P_  clock_i _01342_ \atbs_core_0.spike_memory_0.n2381_o[8]\ _13359_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[446]$_DFFE_PP0P_  clock_i _01343_ \atbs_core_0.spike_memory_0.n2381_o[9]\ _13358_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[447]$_DFFE_PP0P_  clock_i _01344_ \atbs_core_0.spike_memory_0.n2381_o[10]\ _13357_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[448]$_DFFE_PP0P_  clock_i _01345_ \atbs_core_0.spike_memory_0.n2381_o[11]\ _13356_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[449]$_DFFE_PP0P_  clock_i _01346_ \atbs_core_0.spike_memory_0.n2381_o[12]\ _13355_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[44]$_DFFE_PP0P_  clock_i _01347_ \atbs_core_0.spike_memory_0.n2360_o[6]\ _13354_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[450]$_DFFE_PP0P_  clock_i _01348_ \atbs_core_0.spike_memory_0.n2381_o[13]\ _13353_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[451]$_DFFE_PP0P_  clock_i _01349_ \atbs_core_0.spike_memory_0.n2381_o[14]\ _13352_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[452]$_DFFE_PP0P_  clock_i _01350_ \atbs_core_0.spike_memory_0.n2381_o[15]\ _13351_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[453]$_DFFE_PP0P_  clock_i _01351_ \atbs_core_0.spike_memory_0.n2381_o[16]\ _13350_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[454]$_DFFE_PP0P_  clock_i _01352_ \atbs_core_0.spike_memory_0.n2381_o[17]\ _13349_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[455]$_DFFE_PP0P_  clock_i _01353_ \atbs_core_0.spike_memory_0.n2381_o[18]\ _13348_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[456]$_DFFE_PP0P_  clock_i _01354_ \atbs_core_0.spike_memory_0.n2382_o[0]\ _13347_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[457]$_DFFE_PP0P_  clock_i _01355_ \atbs_core_0.spike_memory_0.n2382_o[1]\ _13346_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[458]$_DFFE_PP0P_  clock_i _01356_ \atbs_core_0.spike_memory_0.n2382_o[2]\ _13345_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[459]$_DFFE_PP0P_  clock_i _01357_ \atbs_core_0.spike_memory_0.n2382_o[3]\ _13344_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[45]$_DFFE_PP0P_  clock_i _01358_ \atbs_core_0.spike_memory_0.n2360_o[7]\ _13343_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[460]$_DFFE_PP0P_  clock_i _01359_ \atbs_core_0.spike_memory_0.n2382_o[4]\ _13342_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[461]$_DFFE_PP0P_  clock_i _01360_ \atbs_core_0.spike_memory_0.n2382_o[5]\ _13341_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[462]$_DFFE_PP0P_  clock_i _01361_ \atbs_core_0.spike_memory_0.n2382_o[6]\ _13340_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[463]$_DFFE_PP0P_  clock_i _01362_ \atbs_core_0.spike_memory_0.n2382_o[7]\ _13339_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[464]$_DFFE_PP0P_  clock_i _01363_ \atbs_core_0.spike_memory_0.n2382_o[8]\ _13338_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[465]$_DFFE_PP0P_  clock_i _01364_ \atbs_core_0.spike_memory_0.n2382_o[9]\ _13337_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[466]$_DFFE_PP0P_  clock_i _01365_ \atbs_core_0.spike_memory_0.n2382_o[10]\ _13336_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[467]$_DFFE_PP0P_  clock_i _01366_ \atbs_core_0.spike_memory_0.n2382_o[11]\ _13335_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[468]$_DFFE_PP0P_  clock_i _01367_ \atbs_core_0.spike_memory_0.n2382_o[12]\ _13334_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[469]$_DFFE_PP0P_  clock_i _01368_ \atbs_core_0.spike_memory_0.n2382_o[13]\ _13333_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[46]$_DFFE_PP0P_  clock_i _01369_ \atbs_core_0.spike_memory_0.n2360_o[8]\ _13332_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[470]$_DFFE_PP0P_  clock_i _01370_ \atbs_core_0.spike_memory_0.n2382_o[14]\ _13331_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[471]$_DFFE_PP0P_  clock_i _01371_ \atbs_core_0.spike_memory_0.n2382_o[15]\ _13330_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[472]$_DFFE_PP0P_  clock_i _01372_ \atbs_core_0.spike_memory_0.n2382_o[16]\ _13329_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[473]$_DFFE_PP0P_  clock_i _01373_ \atbs_core_0.spike_memory_0.n2382_o[17]\ _13328_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[474]$_DFFE_PP0P_  clock_i _01374_ \atbs_core_0.spike_memory_0.n2382_o[18]\ _13327_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[475]$_DFFE_PP0P_  clock_i _01375_ \atbs_core_0.spike_memory_0.n2383_o[0]\ _13326_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[476]$_DFFE_PP0P_  clock_i _01376_ \atbs_core_0.spike_memory_0.n2383_o[1]\ _13325_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[477]$_DFFE_PP0P_  clock_i _01377_ \atbs_core_0.spike_memory_0.n2383_o[2]\ _13324_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[478]$_DFFE_PP0P_  clock_i _01378_ \atbs_core_0.spike_memory_0.n2383_o[3]\ _13323_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[479]$_DFFE_PP0P_  clock_i _01379_ \atbs_core_0.spike_memory_0.n2383_o[4]\ _13322_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[47]$_DFFE_PP0P_  clock_i _01380_ \atbs_core_0.spike_memory_0.n2360_o[9]\ _13321_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[480]$_DFFE_PP0P_  clock_i _01381_ \atbs_core_0.spike_memory_0.n2383_o[5]\ _13320_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[481]$_DFFE_PP0P_  clock_i _01382_ \atbs_core_0.spike_memory_0.n2383_o[6]\ _13319_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[482]$_DFFE_PP0P_  clock_i _01383_ \atbs_core_0.spike_memory_0.n2383_o[7]\ _13318_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[483]$_DFFE_PP0P_  clock_i _01384_ \atbs_core_0.spike_memory_0.n2383_o[8]\ _13317_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[484]$_DFFE_PP0P_  clock_i _01385_ \atbs_core_0.spike_memory_0.n2383_o[9]\ _13316_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[485]$_DFFE_PP0P_  clock_i _01386_ \atbs_core_0.spike_memory_0.n2383_o[10]\ _13315_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[486]$_DFFE_PP0P_  clock_i _01387_ \atbs_core_0.spike_memory_0.n2383_o[11]\ _13314_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[487]$_DFFE_PP0P_  clock_i _01388_ \atbs_core_0.spike_memory_0.n2383_o[12]\ _13313_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[488]$_DFFE_PP0P_  clock_i _01389_ \atbs_core_0.spike_memory_0.n2383_o[13]\ _13312_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[489]$_DFFE_PP0P_  clock_i _01390_ \atbs_core_0.spike_memory_0.n2383_o[14]\ _13311_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[48]$_DFFE_PP0P_  clock_i _01391_ \atbs_core_0.spike_memory_0.n2360_o[10]\ _13310_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[490]$_DFFE_PP0P_  clock_i _01392_ \atbs_core_0.spike_memory_0.n2383_o[15]\ _13309_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[491]$_DFFE_PP0P_  clock_i _01393_ \atbs_core_0.spike_memory_0.n2383_o[16]\ _13308_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[492]$_DFFE_PP0P_  clock_i _01394_ \atbs_core_0.spike_memory_0.n2383_o[17]\ _13307_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[493]$_DFFE_PP0P_  clock_i _01395_ \atbs_core_0.spike_memory_0.n2383_o[18]\ _13306_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[494]$_DFFE_PP0P_  clock_i _01396_ \atbs_core_0.spike_memory_0.n2384_o[0]\ _13305_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[495]$_DFFE_PP0P_  clock_i _01397_ \atbs_core_0.spike_memory_0.n2384_o[1]\ _13304_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[496]$_DFFE_PP0P_  clock_i _01398_ \atbs_core_0.spike_memory_0.n2384_o[2]\ _13303_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[497]$_DFFE_PP0P_  clock_i _01399_ \atbs_core_0.spike_memory_0.n2384_o[3]\ _13302_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[498]$_DFFE_PP0P_  clock_i _01400_ \atbs_core_0.spike_memory_0.n2384_o[4]\ _13301_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[499]$_DFFE_PP0P_  clock_i _01401_ \atbs_core_0.spike_memory_0.n2384_o[5]\ _13300_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[49]$_DFFE_PP0P_  clock_i _01402_ \atbs_core_0.spike_memory_0.n2360_o[11]\ _13299_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[4]$_DFFE_PP0P_  clock_i _01403_ \atbs_core_0.spike_memory_0.n2358_o[4]\ _13298_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[500]$_DFFE_PP0P_  clock_i _01404_ \atbs_core_0.spike_memory_0.n2384_o[6]\ _13297_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[501]$_DFFE_PP0P_  clock_i _01405_ \atbs_core_0.spike_memory_0.n2384_o[7]\ _13296_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[502]$_DFFE_PP0P_  clock_i _01406_ \atbs_core_0.spike_memory_0.n2384_o[8]\ _13295_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[503]$_DFFE_PP0P_  clock_i _01407_ \atbs_core_0.spike_memory_0.n2384_o[9]\ _13294_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[504]$_DFFE_PP0P_  clock_i _01408_ \atbs_core_0.spike_memory_0.n2384_o[10]\ _13293_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[505]$_DFFE_PP0P_  clock_i _01409_ \atbs_core_0.spike_memory_0.n2384_o[11]\ _13292_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[506]$_DFFE_PP0P_  clock_i _01410_ \atbs_core_0.spike_memory_0.n2384_o[12]\ _13291_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[507]$_DFFE_PP0P_  clock_i _01411_ \atbs_core_0.spike_memory_0.n2384_o[13]\ _13290_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[508]$_DFFE_PP0P_  clock_i _01412_ \atbs_core_0.spike_memory_0.n2384_o[14]\ _13289_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[509]$_DFFE_PP0P_  clock_i _01413_ \atbs_core_0.spike_memory_0.n2384_o[15]\ _13288_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[50]$_DFFE_PP0P_  clock_i _01414_ \atbs_core_0.spike_memory_0.n2360_o[12]\ _13287_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[510]$_DFFE_PP0P_  clock_i _01415_ \atbs_core_0.spike_memory_0.n2384_o[16]\ _13286_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[511]$_DFFE_PP0P_  clock_i _01416_ \atbs_core_0.spike_memory_0.n2384_o[17]\ _13285_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[512]$_DFFE_PP0P_  clock_i _01417_ \atbs_core_0.spike_memory_0.n2384_o[18]\ _13284_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[513]$_DFFE_PP0P_  clock_i _01418_ \atbs_core_0.spike_memory_0.n2385_o[0]\ _13283_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[514]$_DFFE_PP0P_  clock_i _01419_ \atbs_core_0.spike_memory_0.n2385_o[1]\ _13282_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[515]$_DFFE_PP0P_  clock_i _01420_ \atbs_core_0.spike_memory_0.n2385_o[2]\ _13281_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[516]$_DFFE_PP0P_  clock_i _01421_ \atbs_core_0.spike_memory_0.n2385_o[3]\ _13280_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[517]$_DFFE_PP0P_  clock_i _01422_ \atbs_core_0.spike_memory_0.n2385_o[4]\ _13279_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[518]$_DFFE_PP0P_  clock_i _01423_ \atbs_core_0.spike_memory_0.n2385_o[5]\ _13278_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[519]$_DFFE_PP0P_  clock_i _01424_ \atbs_core_0.spike_memory_0.n2385_o[6]\ _13277_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[51]$_DFFE_PP0P_  clock_i _01425_ \atbs_core_0.spike_memory_0.n2360_o[13]\ _13276_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[520]$_DFFE_PP0P_  clock_i _01426_ \atbs_core_0.spike_memory_0.n2385_o[7]\ _13275_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[521]$_DFFE_PP0P_  clock_i _01427_ \atbs_core_0.spike_memory_0.n2385_o[8]\ _13274_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[522]$_DFFE_PP0P_  clock_i _01428_ \atbs_core_0.spike_memory_0.n2385_o[9]\ _13273_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[523]$_DFFE_PP0P_  clock_i _01429_ \atbs_core_0.spike_memory_0.n2385_o[10]\ _13272_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[524]$_DFFE_PP0P_  clock_i _01430_ \atbs_core_0.spike_memory_0.n2385_o[11]\ _13271_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[525]$_DFFE_PP0P_  clock_i _01431_ \atbs_core_0.spike_memory_0.n2385_o[12]\ _13270_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[526]$_DFFE_PP0P_  clock_i _01432_ \atbs_core_0.spike_memory_0.n2385_o[13]\ _13269_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[527]$_DFFE_PP0P_  clock_i _01433_ \atbs_core_0.spike_memory_0.n2385_o[14]\ _13268_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[528]$_DFFE_PP0P_  clock_i _01434_ \atbs_core_0.spike_memory_0.n2385_o[15]\ _13267_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[529]$_DFFE_PP0P_  clock_i _01435_ \atbs_core_0.spike_memory_0.n2385_o[16]\ _13266_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[52]$_DFFE_PP0P_  clock_i _01436_ \atbs_core_0.spike_memory_0.n2360_o[14]\ _13265_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[530]$_DFFE_PP0P_  clock_i _01437_ \atbs_core_0.spike_memory_0.n2385_o[17]\ _13264_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[531]$_DFFE_PP0P_  clock_i _01438_ \atbs_core_0.spike_memory_0.n2385_o[18]\ _13263_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[532]$_DFFE_PP0P_  clock_i _01439_ \atbs_core_0.spike_memory_0.n2386_o[0]\ _13262_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[533]$_DFFE_PP0P_  clock_i _01440_ \atbs_core_0.spike_memory_0.n2386_o[1]\ _13261_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[534]$_DFFE_PP0P_  clock_i _01441_ \atbs_core_0.spike_memory_0.n2386_o[2]\ _13260_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[535]$_DFFE_PP0P_  clock_i _01442_ \atbs_core_0.spike_memory_0.n2386_o[3]\ _13259_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[536]$_DFFE_PP0P_  clock_i _01443_ \atbs_core_0.spike_memory_0.n2386_o[4]\ _13258_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[537]$_DFFE_PP0P_  clock_i _01444_ \atbs_core_0.spike_memory_0.n2386_o[5]\ _13257_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[538]$_DFFE_PP0P_  clock_i _01445_ \atbs_core_0.spike_memory_0.n2386_o[6]\ _13256_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[539]$_DFFE_PP0P_  clock_i _01446_ \atbs_core_0.spike_memory_0.n2386_o[7]\ _13255_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[53]$_DFFE_PP0P_  clock_i _01447_ \atbs_core_0.spike_memory_0.n2360_o[15]\ _13254_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[540]$_DFFE_PP0P_  clock_i _01448_ \atbs_core_0.spike_memory_0.n2386_o[8]\ _13253_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[541]$_DFFE_PP0P_  clock_i _01449_ \atbs_core_0.spike_memory_0.n2386_o[9]\ _13252_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[542]$_DFFE_PP0P_  clock_i _01450_ \atbs_core_0.spike_memory_0.n2386_o[10]\ _13251_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[543]$_DFFE_PP0P_  clock_i _01451_ \atbs_core_0.spike_memory_0.n2386_o[11]\ _13250_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[544]$_DFFE_PP0P_  clock_i _01452_ \atbs_core_0.spike_memory_0.n2386_o[12]\ _13249_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[545]$_DFFE_PP0P_  clock_i _01453_ \atbs_core_0.spike_memory_0.n2386_o[13]\ _13248_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[546]$_DFFE_PP0P_  clock_i _01454_ \atbs_core_0.spike_memory_0.n2386_o[14]\ _13247_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[547]$_DFFE_PP0P_  clock_i _01455_ \atbs_core_0.spike_memory_0.n2386_o[15]\ _13246_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[548]$_DFFE_PP0P_  clock_i _01456_ \atbs_core_0.spike_memory_0.n2386_o[16]\ _13245_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[549]$_DFFE_PP0P_  clock_i _01457_ \atbs_core_0.spike_memory_0.n2386_o[17]\ _13244_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[54]$_DFFE_PP0P_  clock_i _01458_ \atbs_core_0.spike_memory_0.n2360_o[16]\ _13243_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[550]$_DFFE_PP0P_  clock_i _01459_ \atbs_core_0.spike_memory_0.n2386_o[18]\ _13242_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[551]$_DFFE_PP0P_  clock_i _01460_ \atbs_core_0.spike_memory_0.n2387_o[0]\ _13241_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[552]$_DFFE_PP0P_  clock_i _01461_ \atbs_core_0.spike_memory_0.n2387_o[1]\ _13240_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[553]$_DFFE_PP0P_  clock_i _01462_ \atbs_core_0.spike_memory_0.n2387_o[2]\ _13239_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[554]$_DFFE_PP0P_  clock_i _01463_ \atbs_core_0.spike_memory_0.n2387_o[3]\ _13238_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[555]$_DFFE_PP0P_  clock_i _01464_ \atbs_core_0.spike_memory_0.n2387_o[4]\ _13237_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[556]$_DFFE_PP0P_  clock_i _01465_ \atbs_core_0.spike_memory_0.n2387_o[5]\ _13236_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[557]$_DFFE_PP0P_  clock_i _01466_ \atbs_core_0.spike_memory_0.n2387_o[6]\ _13235_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[558]$_DFFE_PP0P_  clock_i _01467_ \atbs_core_0.spike_memory_0.n2387_o[7]\ _13234_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[559]$_DFFE_PP0P_  clock_i _01468_ \atbs_core_0.spike_memory_0.n2387_o[8]\ _13233_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[55]$_DFFE_PP0P_  clock_i _01469_ \atbs_core_0.spike_memory_0.n2360_o[17]\ _13232_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[560]$_DFFE_PP0P_  clock_i _01470_ \atbs_core_0.spike_memory_0.n2387_o[9]\ _13231_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[561]$_DFFE_PP0P_  clock_i _01471_ \atbs_core_0.spike_memory_0.n2387_o[10]\ _13230_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[562]$_DFFE_PP0P_  clock_i _01472_ \atbs_core_0.spike_memory_0.n2387_o[11]\ _13229_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[563]$_DFFE_PP0P_  clock_i _01473_ \atbs_core_0.spike_memory_0.n2387_o[12]\ _13228_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[564]$_DFFE_PP0P_  clock_i _01474_ \atbs_core_0.spike_memory_0.n2387_o[13]\ _13227_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[565]$_DFFE_PP0P_  clock_i _01475_ \atbs_core_0.spike_memory_0.n2387_o[14]\ _13226_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[566]$_DFFE_PP0P_  clock_i _01476_ \atbs_core_0.spike_memory_0.n2387_o[15]\ _13225_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[567]$_DFFE_PP0P_  clock_i _01477_ \atbs_core_0.spike_memory_0.n2387_o[16]\ _13224_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[568]$_DFFE_PP0P_  clock_i _01478_ \atbs_core_0.spike_memory_0.n2387_o[17]\ _13223_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[569]$_DFFE_PP0P_  clock_i _01479_ \atbs_core_0.spike_memory_0.n2387_o[18]\ _13222_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[56]$_DFFE_PP0P_  clock_i _01480_ \atbs_core_0.spike_memory_0.n2360_o[18]\ _13221_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[570]$_DFFE_PP0P_  clock_i _01481_ \atbs_core_0.spike_memory_0.n2388_o[0]\ _13220_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[571]$_DFFE_PP0P_  clock_i _01482_ \atbs_core_0.spike_memory_0.n2388_o[1]\ _13219_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[572]$_DFFE_PP0P_  clock_i _01483_ \atbs_core_0.spike_memory_0.n2388_o[2]\ _13218_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[573]$_DFFE_PP0P_  clock_i _01484_ \atbs_core_0.spike_memory_0.n2388_o[3]\ _13217_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[574]$_DFFE_PP0P_  clock_i _01485_ \atbs_core_0.spike_memory_0.n2388_o[4]\ _13216_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[575]$_DFFE_PP0P_  clock_i _01486_ \atbs_core_0.spike_memory_0.n2388_o[5]\ _13215_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[576]$_DFFE_PP0P_  clock_i _01487_ \atbs_core_0.spike_memory_0.n2388_o[6]\ _13214_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[577]$_DFFE_PP0P_  clock_i _01488_ \atbs_core_0.spike_memory_0.n2388_o[7]\ _13213_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[578]$_DFFE_PP0P_  clock_i _01489_ \atbs_core_0.spike_memory_0.n2388_o[8]\ _13212_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[579]$_DFFE_PP0P_  clock_i _01490_ \atbs_core_0.spike_memory_0.n2388_o[9]\ _13211_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[57]$_DFFE_PP0P_  clock_i _01491_ \atbs_core_0.spike_memory_0.n2361_o[0]\ _13210_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[580]$_DFFE_PP0P_  clock_i _01492_ \atbs_core_0.spike_memory_0.n2388_o[10]\ _13209_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[581]$_DFFE_PP0P_  clock_i _01493_ \atbs_core_0.spike_memory_0.n2388_o[11]\ _13208_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[582]$_DFFE_PP0P_  clock_i _01494_ \atbs_core_0.spike_memory_0.n2388_o[12]\ _13207_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[583]$_DFFE_PP0P_  clock_i _01495_ \atbs_core_0.spike_memory_0.n2388_o[13]\ _13206_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[584]$_DFFE_PP0P_  clock_i _01496_ \atbs_core_0.spike_memory_0.n2388_o[14]\ _13205_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[585]$_DFFE_PP0P_  clock_i _01497_ \atbs_core_0.spike_memory_0.n2388_o[15]\ _13204_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[586]$_DFFE_PP0P_  clock_i _01498_ \atbs_core_0.spike_memory_0.n2388_o[16]\ _13203_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[587]$_DFFE_PP0P_  clock_i _01499_ \atbs_core_0.spike_memory_0.n2388_o[17]\ _13202_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[588]$_DFFE_PP0P_  clock_i _01500_ \atbs_core_0.spike_memory_0.n2388_o[18]\ _13201_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[589]$_DFFE_PP0P_  clock_i _01501_ \atbs_core_0.spike_memory_0.n2389_o[0]\ _13200_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[58]$_DFFE_PP0P_  clock_i _01502_ \atbs_core_0.spike_memory_0.n2361_o[1]\ _13199_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[590]$_DFFE_PP0P_  clock_i _01503_ \atbs_core_0.spike_memory_0.n2389_o[1]\ _13198_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[591]$_DFFE_PP0P_  clock_i _01504_ \atbs_core_0.spike_memory_0.n2389_o[2]\ _13197_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[592]$_DFFE_PP0P_  clock_i _01505_ \atbs_core_0.spike_memory_0.n2389_o[3]\ _13196_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[593]$_DFFE_PP0P_  clock_i _01506_ \atbs_core_0.spike_memory_0.n2389_o[4]\ _13195_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[594]$_DFFE_PP0P_  clock_i _01507_ \atbs_core_0.spike_memory_0.n2389_o[5]\ _13194_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[595]$_DFFE_PP0P_  clock_i _01508_ \atbs_core_0.spike_memory_0.n2389_o[6]\ _13193_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[596]$_DFFE_PP0P_  clock_i _01509_ \atbs_core_0.spike_memory_0.n2389_o[7]\ _13192_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[597]$_DFFE_PP0P_  clock_i _01510_ \atbs_core_0.spike_memory_0.n2389_o[8]\ _13191_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[598]$_DFFE_PP0P_  clock_i _01511_ \atbs_core_0.spike_memory_0.n2389_o[9]\ _13190_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[599]$_DFFE_PP0P_  clock_i _01512_ \atbs_core_0.spike_memory_0.n2389_o[10]\ _13189_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[59]$_DFFE_PP0P_  clock_i _01513_ \atbs_core_0.spike_memory_0.n2361_o[2]\ _13188_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[5]$_DFFE_PP0P_  clock_i _01514_ \atbs_core_0.spike_memory_0.n2358_o[5]\ _13187_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[600]$_DFFE_PP0P_  clock_i _01515_ \atbs_core_0.spike_memory_0.n2389_o[11]\ _13186_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[601]$_DFFE_PP0P_  clock_i _01516_ \atbs_core_0.spike_memory_0.n2389_o[12]\ _13185_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[602]$_DFFE_PP0P_  clock_i _01517_ \atbs_core_0.spike_memory_0.n2389_o[13]\ _13184_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[603]$_DFFE_PP0P_  clock_i _01518_ \atbs_core_0.spike_memory_0.n2389_o[14]\ _13183_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[604]$_DFFE_PP0P_  clock_i _01519_ \atbs_core_0.spike_memory_0.n2389_o[15]\ _13182_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[605]$_DFFE_PP0P_  clock_i _01520_ \atbs_core_0.spike_memory_0.n2389_o[16]\ _13181_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[606]$_DFFE_PP0P_  clock_i _01521_ \atbs_core_0.spike_memory_0.n2389_o[17]\ _13180_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[607]$_DFFE_PP0P_  clock_i _01522_ \atbs_core_0.spike_memory_0.n2389_o[18]\ _13179_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[608]$_DFFE_PP0P_  clock_i _01523_ \atbs_core_0.spike_memory_0.n2390_o[0]\ _00111_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[609]$_DFFE_PP0P_  clock_i _01524_ \atbs_core_0.spike_memory_0.n2390_o[1]\ _00114_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[60]$_DFFE_PP0P_  clock_i _01525_ \atbs_core_0.spike_memory_0.n2361_o[3]\ _13178_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[610]$_DFFE_PP0P_  clock_i _01526_ \atbs_core_0.spike_memory_0.n2390_o[2]\ _00117_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[611]$_DFFE_PP0P_  clock_i _01527_ \atbs_core_0.spike_memory_0.n2390_o[3]\ _00120_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[612]$_DFFE_PP0P_  clock_i _01528_ \atbs_core_0.spike_memory_0.n2390_o[4]\ _00123_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[613]$_DFFE_PP0P_  clock_i _01529_ \atbs_core_0.spike_memory_0.n2390_o[5]\ _00126_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[614]$_DFFE_PP0P_  clock_i _01530_ \atbs_core_0.spike_memory_0.n2390_o[6]\ _00129_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[615]$_DFFE_PP0P_  clock_i _01531_ \atbs_core_0.spike_memory_0.n2390_o[7]\ _00132_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[616]$_DFFE_PP0P_  clock_i _01532_ \atbs_core_0.spike_memory_0.n2390_o[8]\ _00135_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[617]$_DFFE_PP0P_  clock_i _01533_ \atbs_core_0.spike_memory_0.n2390_o[9]\ _00138_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[618]$_DFFE_PP0P_  clock_i _01534_ \atbs_core_0.spike_memory_0.n2390_o[10]\ _00141_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[619]$_DFFE_PP0P_  clock_i _01535_ \atbs_core_0.spike_memory_0.n2390_o[11]\ _00144_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[61]$_DFFE_PP0P_  clock_i _01536_ \atbs_core_0.spike_memory_0.n2361_o[4]\ _13177_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[620]$_DFFE_PP0P_  clock_i _01537_ \atbs_core_0.spike_memory_0.n2390_o[12]\ _00147_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[621]$_DFFE_PP0P_  clock_i _01538_ \atbs_core_0.spike_memory_0.n2390_o[13]\ _00150_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[622]$_DFFE_PP0P_  clock_i _01539_ \atbs_core_0.spike_memory_0.n2390_o[14]\ _00008_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[623]$_DFFE_PP0P_  clock_i _01540_ \atbs_core_0.spike_memory_0.n2390_o[15]\ _00011_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[624]$_DFFE_PP0P_  clock_i _01541_ \atbs_core_0.spike_memory_0.n2390_o[16]\ _00014_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[625]$_DFFE_PP0P_  clock_i _01542_ \atbs_core_0.spike_memory_0.n2390_o[17]\ _00017_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[626]$_DFFE_PP0P_  clock_i _01543_ \atbs_core_0.spike_memory_0.n2390_o[18]\ _00020_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[627]$_DFFE_PP0P_  clock_i _01544_ \atbs_core_0.spike_memory_0.n2391_o[0]\ _13176_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[628]$_DFFE_PP0P_  clock_i _01545_ \atbs_core_0.spike_memory_0.n2391_o[1]\ _13175_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[629]$_DFFE_PP0P_  clock_i _01546_ \atbs_core_0.spike_memory_0.n2391_o[2]\ _13174_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[62]$_DFFE_PP0P_  clock_i _01547_ \atbs_core_0.spike_memory_0.n2361_o[5]\ _13173_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[630]$_DFFE_PP0P_  clock_i _01548_ \atbs_core_0.spike_memory_0.n2391_o[3]\ _13172_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[631]$_DFFE_PP0P_  clock_i _01549_ \atbs_core_0.spike_memory_0.n2391_o[4]\ _13171_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[632]$_DFFE_PP0P_  clock_i _01550_ \atbs_core_0.spike_memory_0.n2391_o[5]\ _13170_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[633]$_DFFE_PP0P_  clock_i _01551_ \atbs_core_0.spike_memory_0.n2391_o[6]\ _13169_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[634]$_DFFE_PP0P_  clock_i _01552_ \atbs_core_0.spike_memory_0.n2391_o[7]\ _13168_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[635]$_DFFE_PP0P_  clock_i _01553_ \atbs_core_0.spike_memory_0.n2391_o[8]\ _13167_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[636]$_DFFE_PP0P_  clock_i _01554_ \atbs_core_0.spike_memory_0.n2391_o[9]\ _13166_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[637]$_DFFE_PP0P_  clock_i _01555_ \atbs_core_0.spike_memory_0.n2391_o[10]\ _13165_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[638]$_DFFE_PP0P_  clock_i _01556_ \atbs_core_0.spike_memory_0.n2391_o[11]\ _13164_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[639]$_DFFE_PP0P_  clock_i _01557_ \atbs_core_0.spike_memory_0.n2391_o[12]\ _13163_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[63]$_DFFE_PP0P_  clock_i _01558_ \atbs_core_0.spike_memory_0.n2361_o[6]\ _13162_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[640]$_DFFE_PP0P_  clock_i _01559_ \atbs_core_0.spike_memory_0.n2391_o[13]\ _13161_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[641]$_DFFE_PP0P_  clock_i _01560_ \atbs_core_0.spike_memory_0.n2391_o[14]\ _13160_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[642]$_DFFE_PP0P_  clock_i _01561_ \atbs_core_0.spike_memory_0.n2391_o[15]\ _13159_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[643]$_DFFE_PP0P_  clock_i _01562_ \atbs_core_0.spike_memory_0.n2391_o[16]\ _13158_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[644]$_DFFE_PP0P_  clock_i _01563_ \atbs_core_0.spike_memory_0.n2391_o[17]\ _13157_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[645]$_DFFE_PP0P_  clock_i _01564_ \atbs_core_0.spike_memory_0.n2391_o[18]\ _13156_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[646]$_DFFE_PP0P_  clock_i _01565_ \atbs_core_0.spike_memory_0.n2392_o[0]\ _13155_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[647]$_DFFE_PP0P_  clock_i _01566_ \atbs_core_0.spike_memory_0.n2392_o[1]\ _13154_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[648]$_DFFE_PP0P_  clock_i _01567_ \atbs_core_0.spike_memory_0.n2392_o[2]\ _13153_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[649]$_DFFE_PP0P_  clock_i _01568_ \atbs_core_0.spike_memory_0.n2392_o[3]\ _13152_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[64]$_DFFE_PP0P_  clock_i _01569_ \atbs_core_0.spike_memory_0.n2361_o[7]\ _13151_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[650]$_DFFE_PP0P_  clock_i _01570_ \atbs_core_0.spike_memory_0.n2392_o[4]\ _13150_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[651]$_DFFE_PP0P_  clock_i _01571_ \atbs_core_0.spike_memory_0.n2392_o[5]\ _13149_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[652]$_DFFE_PP0P_  clock_i _01572_ \atbs_core_0.spike_memory_0.n2392_o[6]\ _13148_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[653]$_DFFE_PP0P_  clock_i _01573_ \atbs_core_0.spike_memory_0.n2392_o[7]\ _13147_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[654]$_DFFE_PP0P_  clock_i _01574_ \atbs_core_0.spike_memory_0.n2392_o[8]\ _13146_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[655]$_DFFE_PP0P_  clock_i _01575_ \atbs_core_0.spike_memory_0.n2392_o[9]\ _13145_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[656]$_DFFE_PP0P_  clock_i _01576_ \atbs_core_0.spike_memory_0.n2392_o[10]\ _13144_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[657]$_DFFE_PP0P_  clock_i _01577_ \atbs_core_0.spike_memory_0.n2392_o[11]\ _13143_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[658]$_DFFE_PP0P_  clock_i _01578_ \atbs_core_0.spike_memory_0.n2392_o[12]\ _13142_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[659]$_DFFE_PP0P_  clock_i _01579_ \atbs_core_0.spike_memory_0.n2392_o[13]\ _13141_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[65]$_DFFE_PP0P_  clock_i _01580_ \atbs_core_0.spike_memory_0.n2361_o[8]\ _13140_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[660]$_DFFE_PP0P_  clock_i _01581_ \atbs_core_0.spike_memory_0.n2392_o[14]\ _13139_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[661]$_DFFE_PP0P_  clock_i _01582_ \atbs_core_0.spike_memory_0.n2392_o[15]\ _13138_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[662]$_DFFE_PP0P_  clock_i _01583_ \atbs_core_0.spike_memory_0.n2392_o[16]\ _13137_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[663]$_DFFE_PP0P_  clock_i _01584_ \atbs_core_0.spike_memory_0.n2392_o[17]\ _13136_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[664]$_DFFE_PP0P_  clock_i _01585_ \atbs_core_0.spike_memory_0.n2392_o[18]\ _13135_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[665]$_DFFE_PP0P_  clock_i _01586_ \atbs_core_0.spike_memory_0.n2393_o[0]\ _13134_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[666]$_DFFE_PP0P_  clock_i _01587_ \atbs_core_0.spike_memory_0.n2393_o[1]\ _13133_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[667]$_DFFE_PP0P_  clock_i _01588_ \atbs_core_0.spike_memory_0.n2393_o[2]\ _13132_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[668]$_DFFE_PP0P_  clock_i _01589_ \atbs_core_0.spike_memory_0.n2393_o[3]\ _13131_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[669]$_DFFE_PP0P_  clock_i _01590_ \atbs_core_0.spike_memory_0.n2393_o[4]\ _13130_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[66]$_DFFE_PP0P_  clock_i _01591_ \atbs_core_0.spike_memory_0.n2361_o[9]\ _13129_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[670]$_DFFE_PP0P_  clock_i _01592_ \atbs_core_0.spike_memory_0.n2393_o[5]\ _13128_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[671]$_DFFE_PP0P_  clock_i _01593_ \atbs_core_0.spike_memory_0.n2393_o[6]\ _13127_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[672]$_DFFE_PP0P_  clock_i _01594_ \atbs_core_0.spike_memory_0.n2393_o[7]\ _13126_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[673]$_DFFE_PP0P_  clock_i _01595_ \atbs_core_0.spike_memory_0.n2393_o[8]\ _13125_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[674]$_DFFE_PP0P_  clock_i _01596_ \atbs_core_0.spike_memory_0.n2393_o[9]\ _13124_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[675]$_DFFE_PP0P_  clock_i _01597_ \atbs_core_0.spike_memory_0.n2393_o[10]\ _13123_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[676]$_DFFE_PP0P_  clock_i _01598_ \atbs_core_0.spike_memory_0.n2393_o[11]\ _13122_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[677]$_DFFE_PP0P_  clock_i _01599_ \atbs_core_0.spike_memory_0.n2393_o[12]\ _13121_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[678]$_DFFE_PP0P_  clock_i _01600_ \atbs_core_0.spike_memory_0.n2393_o[13]\ _13120_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[679]$_DFFE_PP0P_  clock_i _01601_ \atbs_core_0.spike_memory_0.n2393_o[14]\ _13119_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[67]$_DFFE_PP0P_  clock_i _01602_ \atbs_core_0.spike_memory_0.n2361_o[10]\ _13118_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[680]$_DFFE_PP0P_  clock_i _01603_ \atbs_core_0.spike_memory_0.n2393_o[15]\ _13117_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[681]$_DFFE_PP0P_  clock_i _01604_ \atbs_core_0.spike_memory_0.n2393_o[16]\ _13116_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[682]$_DFFE_PP0P_  clock_i _01605_ \atbs_core_0.spike_memory_0.n2393_o[17]\ _13115_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[683]$_DFFE_PP0P_  clock_i _01606_ \atbs_core_0.spike_memory_0.n2393_o[18]\ _13114_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[684]$_DFFE_PP0P_  clock_i _01607_ \atbs_core_0.spike_memory_0.n2394_o[0]\ _13113_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[685]$_DFFE_PP0P_  clock_i _01608_ \atbs_core_0.spike_memory_0.n2394_o[1]\ _13112_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[686]$_DFFE_PP0P_  clock_i _01609_ \atbs_core_0.spike_memory_0.n2394_o[2]\ _13111_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[687]$_DFFE_PP0P_  clock_i _01610_ \atbs_core_0.spike_memory_0.n2394_o[3]\ _13110_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[688]$_DFFE_PP0P_  clock_i _01611_ \atbs_core_0.spike_memory_0.n2394_o[4]\ _13109_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[689]$_DFFE_PP0P_  clock_i _01612_ \atbs_core_0.spike_memory_0.n2394_o[5]\ _13108_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[68]$_DFFE_PP0P_  clock_i _01613_ \atbs_core_0.spike_memory_0.n2361_o[11]\ _13107_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[690]$_DFFE_PP0P_  clock_i _01614_ \atbs_core_0.spike_memory_0.n2394_o[6]\ _13106_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[691]$_DFFE_PP0P_  clock_i _01615_ \atbs_core_0.spike_memory_0.n2394_o[7]\ _13105_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[692]$_DFFE_PP0P_  clock_i _01616_ \atbs_core_0.spike_memory_0.n2394_o[8]\ _13104_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[693]$_DFFE_PP0P_  clock_i _01617_ \atbs_core_0.spike_memory_0.n2394_o[9]\ _13103_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[694]$_DFFE_PP0P_  clock_i _01618_ \atbs_core_0.spike_memory_0.n2394_o[10]\ _13102_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[695]$_DFFE_PP0P_  clock_i _01619_ \atbs_core_0.spike_memory_0.n2394_o[11]\ _13101_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[696]$_DFFE_PP0P_  clock_i _01620_ \atbs_core_0.spike_memory_0.n2394_o[12]\ _13100_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[697]$_DFFE_PP0P_  clock_i _01621_ \atbs_core_0.spike_memory_0.n2394_o[13]\ _13099_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[698]$_DFFE_PP0P_  clock_i _01622_ \atbs_core_0.spike_memory_0.n2394_o[14]\ _13098_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[699]$_DFFE_PP0P_  clock_i _01623_ \atbs_core_0.spike_memory_0.n2394_o[15]\ _13097_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[69]$_DFFE_PP0P_  clock_i _01624_ \atbs_core_0.spike_memory_0.n2361_o[12]\ _13096_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[6]$_DFFE_PP0P_  clock_i _01625_ \atbs_core_0.spike_memory_0.n2358_o[6]\ _13095_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[700]$_DFFE_PP0P_  clock_i _01626_ \atbs_core_0.spike_memory_0.n2394_o[16]\ _13094_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[701]$_DFFE_PP0P_  clock_i _01627_ \atbs_core_0.spike_memory_0.n2394_o[17]\ _13093_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[702]$_DFFE_PP0P_  clock_i _01628_ \atbs_core_0.spike_memory_0.n2394_o[18]\ _13092_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[703]$_DFFE_PP0P_  clock_i _01629_ \atbs_core_0.spike_memory_0.n2395_o[0]\ _13091_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[704]$_DFFE_PP0P_  clock_i _01630_ \atbs_core_0.spike_memory_0.n2395_o[1]\ _13090_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[705]$_DFFE_PP0P_  clock_i _01631_ \atbs_core_0.spike_memory_0.n2395_o[2]\ _13089_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[706]$_DFFE_PP0P_  clock_i _01632_ \atbs_core_0.spike_memory_0.n2395_o[3]\ _13088_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[707]$_DFFE_PP0P_  clock_i _01633_ \atbs_core_0.spike_memory_0.n2395_o[4]\ _13087_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[708]$_DFFE_PP0P_  clock_i _01634_ \atbs_core_0.spike_memory_0.n2395_o[5]\ _13086_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[709]$_DFFE_PP0P_  clock_i _01635_ \atbs_core_0.spike_memory_0.n2395_o[6]\ _13085_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[70]$_DFFE_PP0P_  clock_i _01636_ \atbs_core_0.spike_memory_0.n2361_o[13]\ _13084_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[710]$_DFFE_PP0P_  clock_i _01637_ \atbs_core_0.spike_memory_0.n2395_o[7]\ _13083_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[711]$_DFFE_PP0P_  clock_i _01638_ \atbs_core_0.spike_memory_0.n2395_o[8]\ _13082_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[712]$_DFFE_PP0P_  clock_i _01639_ \atbs_core_0.spike_memory_0.n2395_o[9]\ _13081_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[713]$_DFFE_PP0P_  clock_i _01640_ \atbs_core_0.spike_memory_0.n2395_o[10]\ _13080_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[714]$_DFFE_PP0P_  clock_i _01641_ \atbs_core_0.spike_memory_0.n2395_o[11]\ _13079_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[715]$_DFFE_PP0P_  clock_i _01642_ \atbs_core_0.spike_memory_0.n2395_o[12]\ _13078_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[716]$_DFFE_PP0P_  clock_i _01643_ \atbs_core_0.spike_memory_0.n2395_o[13]\ _13077_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[717]$_DFFE_PP0P_  clock_i _01644_ \atbs_core_0.spike_memory_0.n2395_o[14]\ _13076_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[718]$_DFFE_PP0P_  clock_i _01645_ \atbs_core_0.spike_memory_0.n2395_o[15]\ _13075_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[719]$_DFFE_PP0P_  clock_i _01646_ \atbs_core_0.spike_memory_0.n2395_o[16]\ _13074_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[71]$_DFFE_PP0P_  clock_i _01647_ \atbs_core_0.spike_memory_0.n2361_o[14]\ _13073_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[720]$_DFFE_PP0P_  clock_i _01648_ \atbs_core_0.spike_memory_0.n2395_o[17]\ _13072_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[721]$_DFFE_PP0P_  clock_i _01649_ \atbs_core_0.spike_memory_0.n2395_o[18]\ _13071_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[722]$_DFFE_PP0P_  clock_i _01650_ \atbs_core_0.spike_memory_0.n2396_o[0]\ _13070_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[723]$_DFFE_PP0P_  clock_i _01651_ \atbs_core_0.spike_memory_0.n2396_o[1]\ _13069_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[724]$_DFFE_PP0P_  clock_i _01652_ \atbs_core_0.spike_memory_0.n2396_o[2]\ _13068_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[725]$_DFFE_PP0P_  clock_i _01653_ \atbs_core_0.spike_memory_0.n2396_o[3]\ _13067_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[726]$_DFFE_PP0P_  clock_i _01654_ \atbs_core_0.spike_memory_0.n2396_o[4]\ _13066_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[727]$_DFFE_PP0P_  clock_i _01655_ \atbs_core_0.spike_memory_0.n2396_o[5]\ _13065_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[728]$_DFFE_PP0P_  clock_i _01656_ \atbs_core_0.spike_memory_0.n2396_o[6]\ _13064_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[729]$_DFFE_PP0P_  clock_i _01657_ \atbs_core_0.spike_memory_0.n2396_o[7]\ _13063_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[72]$_DFFE_PP0P_  clock_i _01658_ \atbs_core_0.spike_memory_0.n2361_o[15]\ _13062_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[730]$_DFFE_PP0P_  clock_i _01659_ \atbs_core_0.spike_memory_0.n2396_o[8]\ _13061_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[731]$_DFFE_PP0P_  clock_i _01660_ \atbs_core_0.spike_memory_0.n2396_o[9]\ _13060_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[732]$_DFFE_PP0P_  clock_i _01661_ \atbs_core_0.spike_memory_0.n2396_o[10]\ _13059_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[733]$_DFFE_PP0P_  clock_i _01662_ \atbs_core_0.spike_memory_0.n2396_o[11]\ _13058_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[734]$_DFFE_PP0P_  clock_i _01663_ \atbs_core_0.spike_memory_0.n2396_o[12]\ _13057_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[735]$_DFFE_PP0P_  clock_i _01664_ \atbs_core_0.spike_memory_0.n2396_o[13]\ _13056_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[736]$_DFFE_PP0P_  clock_i _01665_ \atbs_core_0.spike_memory_0.n2396_o[14]\ _13055_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[737]$_DFFE_PP0P_  clock_i _01666_ \atbs_core_0.spike_memory_0.n2396_o[15]\ _13054_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[738]$_DFFE_PP0P_  clock_i _01667_ \atbs_core_0.spike_memory_0.n2396_o[16]\ _13053_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[739]$_DFFE_PP0P_  clock_i _01668_ \atbs_core_0.spike_memory_0.n2396_o[17]\ _13052_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[73]$_DFFE_PP0P_  clock_i _01669_ \atbs_core_0.spike_memory_0.n2361_o[16]\ _13051_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[740]$_DFFE_PP0P_  clock_i _01670_ \atbs_core_0.spike_memory_0.n2396_o[18]\ _13050_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[741]$_DFFE_PP0P_  clock_i _01671_ \atbs_core_0.spike_memory_0.n2397_o[0]\ _13049_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[742]$_DFFE_PP0P_  clock_i _01672_ \atbs_core_0.spike_memory_0.n2397_o[1]\ _13048_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[743]$_DFFE_PP0P_  clock_i _01673_ \atbs_core_0.spike_memory_0.n2397_o[2]\ _13047_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[744]$_DFFE_PP0P_  clock_i _01674_ \atbs_core_0.spike_memory_0.n2397_o[3]\ _13046_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[745]$_DFFE_PP0P_  clock_i _01675_ \atbs_core_0.spike_memory_0.n2397_o[4]\ _13045_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[746]$_DFFE_PP0P_  clock_i _01676_ \atbs_core_0.spike_memory_0.n2397_o[5]\ _13044_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[747]$_DFFE_PP0P_  clock_i _01677_ \atbs_core_0.spike_memory_0.n2397_o[6]\ _13043_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[748]$_DFFE_PP0P_  clock_i _01678_ \atbs_core_0.spike_memory_0.n2397_o[7]\ _13042_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[749]$_DFFE_PP0P_  clock_i _01679_ \atbs_core_0.spike_memory_0.n2397_o[8]\ _13041_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[74]$_DFFE_PP0P_  clock_i _01680_ \atbs_core_0.spike_memory_0.n2361_o[17]\ _13040_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[750]$_DFFE_PP0P_  clock_i _01681_ \atbs_core_0.spike_memory_0.n2397_o[9]\ _13039_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[751]$_DFFE_PP0P_  clock_i _01682_ \atbs_core_0.spike_memory_0.n2397_o[10]\ _13038_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[752]$_DFFE_PP0P_  clock_i _01683_ \atbs_core_0.spike_memory_0.n2397_o[11]\ _13037_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[753]$_DFFE_PP0P_  clock_i _01684_ \atbs_core_0.spike_memory_0.n2397_o[12]\ _13036_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[754]$_DFFE_PP0P_  clock_i _01685_ \atbs_core_0.spike_memory_0.n2397_o[13]\ _13035_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[755]$_DFFE_PP0P_  clock_i _01686_ \atbs_core_0.spike_memory_0.n2397_o[14]\ _13034_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[756]$_DFFE_PP0P_  clock_i _01687_ \atbs_core_0.spike_memory_0.n2397_o[15]\ _13033_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[757]$_DFFE_PP0P_  clock_i _01688_ \atbs_core_0.spike_memory_0.n2397_o[16]\ _13032_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[758]$_DFFE_PP0P_  clock_i _01689_ \atbs_core_0.spike_memory_0.n2397_o[17]\ _13031_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[759]$_DFFE_PP0P_  clock_i _01690_ \atbs_core_0.spike_memory_0.n2397_o[18]\ _13030_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[75]$_DFFE_PP0P_  clock_i _01691_ \atbs_core_0.spike_memory_0.n2361_o[18]\ _13029_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[760]$_DFFE_PP0P_  clock_i _01692_ \atbs_core_0.spike_memory_0.n2398_o[0]\ _13028_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[761]$_DFFE_PP0P_  clock_i _01693_ \atbs_core_0.spike_memory_0.n2398_o[1]\ _13027_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[762]$_DFFE_PP0P_  clock_i _01694_ \atbs_core_0.spike_memory_0.n2398_o[2]\ _13026_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[763]$_DFFE_PP0P_  clock_i _01695_ \atbs_core_0.spike_memory_0.n2398_o[3]\ _13025_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[764]$_DFFE_PP0P_  clock_i _01696_ \atbs_core_0.spike_memory_0.n2398_o[4]\ _13024_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[765]$_DFFE_PP0P_  clock_i _01697_ \atbs_core_0.spike_memory_0.n2398_o[5]\ _13023_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[766]$_DFFE_PP0P_  clock_i _01698_ \atbs_core_0.spike_memory_0.n2398_o[6]\ _13022_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[767]$_DFFE_PP0P_  clock_i _01699_ \atbs_core_0.spike_memory_0.n2398_o[7]\ _13021_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[768]$_DFFE_PP0P_  clock_i _01700_ \atbs_core_0.spike_memory_0.n2398_o[8]\ _13020_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[769]$_DFFE_PP0P_  clock_i _01701_ \atbs_core_0.spike_memory_0.n2398_o[9]\ _13019_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[76]$_DFFE_PP0P_  clock_i _01702_ \atbs_core_0.spike_memory_0.n2362_o[0]\ _13018_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[770]$_DFFE_PP0P_  clock_i _01703_ \atbs_core_0.spike_memory_0.n2398_o[10]\ _13017_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[771]$_DFFE_PP0P_  clock_i _01704_ \atbs_core_0.spike_memory_0.n2398_o[11]\ _13016_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[772]$_DFFE_PP0P_  clock_i _01705_ \atbs_core_0.spike_memory_0.n2398_o[12]\ _13015_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[773]$_DFFE_PP0P_  clock_i _01706_ \atbs_core_0.spike_memory_0.n2398_o[13]\ _13014_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[774]$_DFFE_PP0P_  clock_i _01707_ \atbs_core_0.spike_memory_0.n2398_o[14]\ _13013_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[775]$_DFFE_PP0P_  clock_i _01708_ \atbs_core_0.spike_memory_0.n2398_o[15]\ _13012_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[776]$_DFFE_PP0P_  clock_i _01709_ \atbs_core_0.spike_memory_0.n2398_o[16]\ _13011_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[777]$_DFFE_PP0P_  clock_i _01710_ \atbs_core_0.spike_memory_0.n2398_o[17]\ _13010_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[778]$_DFFE_PP0P_  clock_i _01711_ \atbs_core_0.spike_memory_0.n2398_o[18]\ _13009_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[779]$_DFFE_PP0P_  clock_i _01712_ \atbs_core_0.spike_memory_0.n2399_o[0]\ _13008_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[77]$_DFFE_PP0P_  clock_i _01713_ \atbs_core_0.spike_memory_0.n2362_o[1]\ _13007_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[780]$_DFFE_PP0P_  clock_i _01714_ \atbs_core_0.spike_memory_0.n2399_o[1]\ _13006_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[781]$_DFFE_PP0P_  clock_i _01715_ \atbs_core_0.spike_memory_0.n2399_o[2]\ _13005_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[782]$_DFFE_PP0P_  clock_i _01716_ \atbs_core_0.spike_memory_0.n2399_o[3]\ _13004_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[783]$_DFFE_PP0P_  clock_i _01717_ \atbs_core_0.spike_memory_0.n2399_o[4]\ _13003_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[784]$_DFFE_PP0P_  clock_i _01718_ \atbs_core_0.spike_memory_0.n2399_o[5]\ _13002_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[785]$_DFFE_PP0P_  clock_i _01719_ \atbs_core_0.spike_memory_0.n2399_o[6]\ _13001_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[786]$_DFFE_PP0P_  clock_i _01720_ \atbs_core_0.spike_memory_0.n2399_o[7]\ _13000_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[787]$_DFFE_PP0P_  clock_i _01721_ \atbs_core_0.spike_memory_0.n2399_o[8]\ _12999_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[788]$_DFFE_PP0P_  clock_i _01722_ \atbs_core_0.spike_memory_0.n2399_o[9]\ _12998_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[789]$_DFFE_PP0P_  clock_i _01723_ \atbs_core_0.spike_memory_0.n2399_o[10]\ _12997_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[78]$_DFFE_PP0P_  clock_i _01724_ \atbs_core_0.spike_memory_0.n2362_o[2]\ _12996_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[790]$_DFFE_PP0P_  clock_i _01725_ \atbs_core_0.spike_memory_0.n2399_o[11]\ _12995_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[791]$_DFFE_PP0P_  clock_i _01726_ \atbs_core_0.spike_memory_0.n2399_o[12]\ _12994_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[792]$_DFFE_PP0P_  clock_i _01727_ \atbs_core_0.spike_memory_0.n2399_o[13]\ _12993_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[793]$_DFFE_PP0P_  clock_i _01728_ \atbs_core_0.spike_memory_0.n2399_o[14]\ _12992_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[794]$_DFFE_PP0P_  clock_i _01729_ \atbs_core_0.spike_memory_0.n2399_o[15]\ _12991_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[795]$_DFFE_PP0P_  clock_i _01730_ \atbs_core_0.spike_memory_0.n2399_o[16]\ _12990_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[796]$_DFFE_PP0P_  clock_i _01731_ \atbs_core_0.spike_memory_0.n2399_o[17]\ _12989_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[797]$_DFFE_PP0P_  clock_i _01732_ \atbs_core_0.spike_memory_0.n2399_o[18]\ _12988_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[798]$_DFFE_PP0P_  clock_i _01733_ \atbs_core_0.spike_memory_0.n2400_o[0]\ _12987_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[799]$_DFFE_PP0P_  clock_i _01734_ \atbs_core_0.spike_memory_0.n2400_o[1]\ _12986_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[79]$_DFFE_PP0P_  clock_i _01735_ \atbs_core_0.spike_memory_0.n2362_o[3]\ _12985_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[7]$_DFFE_PP0P_  clock_i _01736_ \atbs_core_0.spike_memory_0.n2358_o[7]\ _12984_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[800]$_DFFE_PP0P_  clock_i _01737_ \atbs_core_0.spike_memory_0.n2400_o[2]\ _12983_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[801]$_DFFE_PP0P_  clock_i _01738_ \atbs_core_0.spike_memory_0.n2400_o[3]\ _12982_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[802]$_DFFE_PP0P_  clock_i _01739_ \atbs_core_0.spike_memory_0.n2400_o[4]\ _12981_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[803]$_DFFE_PP0P_  clock_i _01740_ \atbs_core_0.spike_memory_0.n2400_o[5]\ _12980_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[804]$_DFFE_PP0P_  clock_i _01741_ \atbs_core_0.spike_memory_0.n2400_o[6]\ _12979_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[805]$_DFFE_PP0P_  clock_i _01742_ \atbs_core_0.spike_memory_0.n2400_o[7]\ _12978_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[806]$_DFFE_PP0P_  clock_i _01743_ \atbs_core_0.spike_memory_0.n2400_o[8]\ _12977_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[807]$_DFFE_PP0P_  clock_i _01744_ \atbs_core_0.spike_memory_0.n2400_o[9]\ _12976_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[808]$_DFFE_PP0P_  clock_i _01745_ \atbs_core_0.spike_memory_0.n2400_o[10]\ _12975_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[809]$_DFFE_PP0P_  clock_i _01746_ \atbs_core_0.spike_memory_0.n2400_o[11]\ _12974_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[80]$_DFFE_PP0P_  clock_i _01747_ \atbs_core_0.spike_memory_0.n2362_o[4]\ _12973_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[810]$_DFFE_PP0P_  clock_i _01748_ \atbs_core_0.spike_memory_0.n2400_o[12]\ _12972_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[811]$_DFFE_PP0P_  clock_i _01749_ \atbs_core_0.spike_memory_0.n2400_o[13]\ _12971_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[812]$_DFFE_PP0P_  clock_i _01750_ \atbs_core_0.spike_memory_0.n2400_o[14]\ _12970_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[813]$_DFFE_PP0P_  clock_i _01751_ \atbs_core_0.spike_memory_0.n2400_o[15]\ _12969_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[814]$_DFFE_PP0P_  clock_i _01752_ \atbs_core_0.spike_memory_0.n2400_o[16]\ _12968_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[815]$_DFFE_PP0P_  clock_i _01753_ \atbs_core_0.spike_memory_0.n2400_o[17]\ _12967_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[816]$_DFFE_PP0P_  clock_i _01754_ \atbs_core_0.spike_memory_0.n2400_o[18]\ _12966_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[817]$_DFFE_PP0P_  clock_i _01755_ \atbs_core_0.spike_memory_0.n2401_o[0]\ _12965_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[818]$_DFFE_PP0P_  clock_i _01756_ \atbs_core_0.spike_memory_0.n2401_o[1]\ _12964_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[819]$_DFFE_PP0P_  clock_i _01757_ \atbs_core_0.spike_memory_0.n2401_o[2]\ _12963_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[81]$_DFFE_PP0P_  clock_i _01758_ \atbs_core_0.spike_memory_0.n2362_o[5]\ _12962_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[820]$_DFFE_PP0P_  clock_i _01759_ \atbs_core_0.spike_memory_0.n2401_o[3]\ _12961_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[821]$_DFFE_PP0P_  clock_i _01760_ \atbs_core_0.spike_memory_0.n2401_o[4]\ _12960_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[822]$_DFFE_PP0P_  clock_i _01761_ \atbs_core_0.spike_memory_0.n2401_o[5]\ _12959_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[823]$_DFFE_PP0P_  clock_i _01762_ \atbs_core_0.spike_memory_0.n2401_o[6]\ _12958_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[824]$_DFFE_PP0P_  clock_i _01763_ \atbs_core_0.spike_memory_0.n2401_o[7]\ _12957_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[825]$_DFFE_PP0P_  clock_i _01764_ \atbs_core_0.spike_memory_0.n2401_o[8]\ _12956_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[826]$_DFFE_PP0P_  clock_i _01765_ \atbs_core_0.spike_memory_0.n2401_o[9]\ _12955_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[827]$_DFFE_PP0P_  clock_i _01766_ \atbs_core_0.spike_memory_0.n2401_o[10]\ _12954_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[828]$_DFFE_PP0P_  clock_i _01767_ \atbs_core_0.spike_memory_0.n2401_o[11]\ _12953_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[829]$_DFFE_PP0P_  clock_i _01768_ \atbs_core_0.spike_memory_0.n2401_o[12]\ _12952_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[82]$_DFFE_PP0P_  clock_i _01769_ \atbs_core_0.spike_memory_0.n2362_o[6]\ _12951_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[830]$_DFFE_PP0P_  clock_i _01770_ \atbs_core_0.spike_memory_0.n2401_o[13]\ _12950_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[831]$_DFFE_PP0P_  clock_i _01771_ \atbs_core_0.spike_memory_0.n2401_o[14]\ _12949_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[832]$_DFFE_PP0P_  clock_i _01772_ \atbs_core_0.spike_memory_0.n2401_o[15]\ _12948_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[833]$_DFFE_PP0P_  clock_i _01773_ \atbs_core_0.spike_memory_0.n2401_o[16]\ _12947_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[834]$_DFFE_PP0P_  clock_i _01774_ \atbs_core_0.spike_memory_0.n2401_o[17]\ _12946_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[835]$_DFFE_PP0P_  clock_i _01775_ \atbs_core_0.spike_memory_0.n2401_o[18]\ _12945_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[836]$_DFFE_PP0P_  clock_i _01776_ \atbs_core_0.spike_memory_0.n2402_o[0]\ _12944_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[837]$_DFFE_PP0P_  clock_i _01777_ \atbs_core_0.spike_memory_0.n2402_o[1]\ _12943_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[838]$_DFFE_PP0P_  clock_i _01778_ \atbs_core_0.spike_memory_0.n2402_o[2]\ _12942_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[839]$_DFFE_PP0P_  clock_i _01779_ \atbs_core_0.spike_memory_0.n2402_o[3]\ _12941_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[83]$_DFFE_PP0P_  clock_i _01780_ \atbs_core_0.spike_memory_0.n2362_o[7]\ _12940_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[840]$_DFFE_PP0P_  clock_i _01781_ \atbs_core_0.spike_memory_0.n2402_o[4]\ _12939_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[841]$_DFFE_PP0P_  clock_i _01782_ \atbs_core_0.spike_memory_0.n2402_o[5]\ _12938_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[842]$_DFFE_PP0P_  clock_i _01783_ \atbs_core_0.spike_memory_0.n2402_o[6]\ _12937_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[843]$_DFFE_PP0P_  clock_i _01784_ \atbs_core_0.spike_memory_0.n2402_o[7]\ _12936_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[844]$_DFFE_PP0P_  clock_i _01785_ \atbs_core_0.spike_memory_0.n2402_o[8]\ _12935_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[845]$_DFFE_PP0P_  clock_i _01786_ \atbs_core_0.spike_memory_0.n2402_o[9]\ _12934_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[846]$_DFFE_PP0P_  clock_i _01787_ \atbs_core_0.spike_memory_0.n2402_o[10]\ _12933_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[847]$_DFFE_PP0P_  clock_i _01788_ \atbs_core_0.spike_memory_0.n2402_o[11]\ _12932_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[848]$_DFFE_PP0P_  clock_i _01789_ \atbs_core_0.spike_memory_0.n2402_o[12]\ _12931_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[849]$_DFFE_PP0P_  clock_i _01790_ \atbs_core_0.spike_memory_0.n2402_o[13]\ _12930_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[84]$_DFFE_PP0P_  clock_i _01791_ \atbs_core_0.spike_memory_0.n2362_o[8]\ _12929_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[850]$_DFFE_PP0P_  clock_i _01792_ \atbs_core_0.spike_memory_0.n2402_o[14]\ _12928_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[851]$_DFFE_PP0P_  clock_i _01793_ \atbs_core_0.spike_memory_0.n2402_o[15]\ _12927_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[852]$_DFFE_PP0P_  clock_i _01794_ \atbs_core_0.spike_memory_0.n2402_o[16]\ _12926_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[853]$_DFFE_PP0P_  clock_i _01795_ \atbs_core_0.spike_memory_0.n2402_o[17]\ _12925_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[854]$_DFFE_PP0P_  clock_i _01796_ \atbs_core_0.spike_memory_0.n2402_o[18]\ _12924_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[855]$_DFFE_PP0P_  clock_i _01797_ \atbs_core_0.spike_memory_0.n2403_o[0]\ _12923_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[856]$_DFFE_PP0P_  clock_i _01798_ \atbs_core_0.spike_memory_0.n2403_o[1]\ _12922_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[857]$_DFFE_PP0P_  clock_i _01799_ \atbs_core_0.spike_memory_0.n2403_o[2]\ _12921_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[858]$_DFFE_PP0P_  clock_i _01800_ \atbs_core_0.spike_memory_0.n2403_o[3]\ _12920_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[859]$_DFFE_PP0P_  clock_i _01801_ \atbs_core_0.spike_memory_0.n2403_o[4]\ _12919_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[85]$_DFFE_PP0P_  clock_i _01802_ \atbs_core_0.spike_memory_0.n2362_o[9]\ _12918_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[860]$_DFFE_PP0P_  clock_i _01803_ \atbs_core_0.spike_memory_0.n2403_o[5]\ _12917_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[861]$_DFFE_PP0P_  clock_i _01804_ \atbs_core_0.spike_memory_0.n2403_o[6]\ _12916_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[862]$_DFFE_PP0P_  clock_i _01805_ \atbs_core_0.spike_memory_0.n2403_o[7]\ _12915_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[863]$_DFFE_PP0P_  clock_i _01806_ \atbs_core_0.spike_memory_0.n2403_o[8]\ _12914_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[864]$_DFFE_PP0P_  clock_i _01807_ \atbs_core_0.spike_memory_0.n2403_o[9]\ _12913_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[865]$_DFFE_PP0P_  clock_i _01808_ \atbs_core_0.spike_memory_0.n2403_o[10]\ _12912_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[866]$_DFFE_PP0P_  clock_i _01809_ \atbs_core_0.spike_memory_0.n2403_o[11]\ _12911_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[867]$_DFFE_PP0P_  clock_i _01810_ \atbs_core_0.spike_memory_0.n2403_o[12]\ _12910_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[868]$_DFFE_PP0P_  clock_i _01811_ \atbs_core_0.spike_memory_0.n2403_o[13]\ _12909_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[869]$_DFFE_PP0P_  clock_i _01812_ \atbs_core_0.spike_memory_0.n2403_o[14]\ _12908_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[86]$_DFFE_PP0P_  clock_i _01813_ \atbs_core_0.spike_memory_0.n2362_o[10]\ _12907_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[870]$_DFFE_PP0P_  clock_i _01814_ \atbs_core_0.spike_memory_0.n2403_o[15]\ _12906_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[871]$_DFFE_PP0P_  clock_i _01815_ \atbs_core_0.spike_memory_0.n2403_o[16]\ _12905_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[872]$_DFFE_PP0P_  clock_i _01816_ \atbs_core_0.spike_memory_0.n2403_o[17]\ _12904_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[873]$_DFFE_PP0P_  clock_i _01817_ \atbs_core_0.spike_memory_0.n2403_o[18]\ _12903_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[874]$_DFFE_PP0P_  clock_i _01818_ \atbs_core_0.spike_memory_0.n2404_o[0]\ _12902_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[875]$_DFFE_PP0P_  clock_i _01819_ \atbs_core_0.spike_memory_0.n2404_o[1]\ _12901_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[876]$_DFFE_PP0P_  clock_i _01820_ \atbs_core_0.spike_memory_0.n2404_o[2]\ _12900_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[877]$_DFFE_PP0P_  clock_i _01821_ \atbs_core_0.spike_memory_0.n2404_o[3]\ _12899_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[878]$_DFFE_PP0P_  clock_i _01822_ \atbs_core_0.spike_memory_0.n2404_o[4]\ _12898_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[879]$_DFFE_PP0P_  clock_i _01823_ \atbs_core_0.spike_memory_0.n2404_o[5]\ _12897_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[87]$_DFFE_PP0P_  clock_i _01824_ \atbs_core_0.spike_memory_0.n2362_o[11]\ _12896_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[880]$_DFFE_PP0P_  clock_i _01825_ \atbs_core_0.spike_memory_0.n2404_o[6]\ _12895_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[881]$_DFFE_PP0P_  clock_i _01826_ \atbs_core_0.spike_memory_0.n2404_o[7]\ _12894_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[882]$_DFFE_PP0P_  clock_i _01827_ \atbs_core_0.spike_memory_0.n2404_o[8]\ _12893_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[883]$_DFFE_PP0P_  clock_i _01828_ \atbs_core_0.spike_memory_0.n2404_o[9]\ _12892_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[884]$_DFFE_PP0P_  clock_i _01829_ \atbs_core_0.spike_memory_0.n2404_o[10]\ _12891_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[885]$_DFFE_PP0P_  clock_i _01830_ \atbs_core_0.spike_memory_0.n2404_o[11]\ _12890_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[886]$_DFFE_PP0P_  clock_i _01831_ \atbs_core_0.spike_memory_0.n2404_o[12]\ _12889_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[887]$_DFFE_PP0P_  clock_i _01832_ \atbs_core_0.spike_memory_0.n2404_o[13]\ _12888_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[888]$_DFFE_PP0P_  clock_i _01833_ \atbs_core_0.spike_memory_0.n2404_o[14]\ _12887_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[889]$_DFFE_PP0P_  clock_i _01834_ \atbs_core_0.spike_memory_0.n2404_o[15]\ _12886_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[88]$_DFFE_PP0P_  clock_i _01835_ \atbs_core_0.spike_memory_0.n2362_o[12]\ _12885_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[890]$_DFFE_PP0P_  clock_i _01836_ \atbs_core_0.spike_memory_0.n2404_o[16]\ _12884_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[891]$_DFFE_PP0P_  clock_i _01837_ \atbs_core_0.spike_memory_0.n2404_o[17]\ _12883_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[892]$_DFFE_PP0P_  clock_i _01838_ \atbs_core_0.spike_memory_0.n2404_o[18]\ _12882_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[893]$_DFFE_PP0P_  clock_i _01839_ \atbs_core_0.spike_memory_0.n2405_o[0]\ _12881_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[894]$_DFFE_PP0P_  clock_i _01840_ \atbs_core_0.spike_memory_0.n2405_o[1]\ _12880_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[895]$_DFFE_PP0P_  clock_i _01841_ \atbs_core_0.spike_memory_0.n2405_o[2]\ _12879_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[896]$_DFFE_PP0P_  clock_i _01842_ \atbs_core_0.spike_memory_0.n2405_o[3]\ _12878_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[897]$_DFFE_PP0P_  clock_i _01843_ \atbs_core_0.spike_memory_0.n2405_o[4]\ _12877_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[898]$_DFFE_PP0P_  clock_i _01844_ \atbs_core_0.spike_memory_0.n2405_o[5]\ _12876_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[899]$_DFFE_PP0P_  clock_i _01845_ \atbs_core_0.spike_memory_0.n2405_o[6]\ _12875_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[89]$_DFFE_PP0P_  clock_i _01846_ \atbs_core_0.spike_memory_0.n2362_o[13]\ _12874_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[8]$_DFFE_PP0P_  clock_i _01847_ \atbs_core_0.spike_memory_0.n2358_o[8]\ _12873_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[900]$_DFFE_PP0P_  clock_i _01848_ \atbs_core_0.spike_memory_0.n2405_o[7]\ _12872_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[901]$_DFFE_PP0P_  clock_i _01849_ \atbs_core_0.spike_memory_0.n2405_o[8]\ _12871_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[902]$_DFFE_PP0P_  clock_i _01850_ \atbs_core_0.spike_memory_0.n2405_o[9]\ _12870_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[903]$_DFFE_PP0P_  clock_i _01851_ \atbs_core_0.spike_memory_0.n2405_o[10]\ _12869_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[904]$_DFFE_PP0P_  clock_i _01852_ \atbs_core_0.spike_memory_0.n2405_o[11]\ _12868_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[905]$_DFFE_PP0P_  clock_i _01853_ \atbs_core_0.spike_memory_0.n2405_o[12]\ _12867_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[906]$_DFFE_PP0P_  clock_i _01854_ \atbs_core_0.spike_memory_0.n2405_o[13]\ _12866_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[907]$_DFFE_PP0P_  clock_i _01855_ \atbs_core_0.spike_memory_0.n2405_o[14]\ _12865_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[908]$_DFFE_PP0P_  clock_i _01856_ \atbs_core_0.spike_memory_0.n2405_o[15]\ _12864_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[909]$_DFFE_PP0P_  clock_i _01857_ \atbs_core_0.spike_memory_0.n2405_o[16]\ _12863_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[90]$_DFFE_PP0P_  clock_i _01858_ \atbs_core_0.spike_memory_0.n2362_o[14]\ _12862_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[910]$_DFFE_PP0P_  clock_i _01859_ \atbs_core_0.spike_memory_0.n2405_o[17]\ _12861_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[911]$_DFFE_PP0P_  clock_i _01860_ \atbs_core_0.spike_memory_0.n2405_o[18]\ _12860_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[912]$_DFFE_PP0P_  clock_i _01861_ \atbs_core_0.spike_memory_0.n2406_o[0]\ _00110_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[913]$_DFFE_PP0P_  clock_i _01862_ \atbs_core_0.spike_memory_0.n2406_o[1]\ _00113_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[914]$_DFFE_PP0P_  clock_i _01863_ \atbs_core_0.spike_memory_0.n2406_o[2]\ _00116_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[915]$_DFFE_PP0P_  clock_i _01864_ \atbs_core_0.spike_memory_0.n2406_o[3]\ _00119_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[916]$_DFFE_PP0P_  clock_i _01865_ \atbs_core_0.spike_memory_0.n2406_o[4]\ _00122_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[917]$_DFFE_PP0P_  clock_i _01866_ \atbs_core_0.spike_memory_0.n2406_o[5]\ _00125_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[918]$_DFFE_PP0P_  clock_i _01867_ \atbs_core_0.spike_memory_0.n2406_o[6]\ _00128_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[919]$_DFFE_PP0P_  clock_i _01868_ \atbs_core_0.spike_memory_0.n2406_o[7]\ _00131_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[91]$_DFFE_PP0P_  clock_i _01869_ \atbs_core_0.spike_memory_0.n2362_o[15]\ _12859_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[920]$_DFFE_PP0P_  clock_i _01870_ \atbs_core_0.spike_memory_0.n2406_o[8]\ _00134_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[921]$_DFFE_PP0P_  clock_i _01871_ \atbs_core_0.spike_memory_0.n2406_o[9]\ _00137_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[922]$_DFFE_PP0P_  clock_i _01872_ \atbs_core_0.spike_memory_0.n2406_o[10]\ _00140_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[923]$_DFFE_PP0P_  clock_i _01873_ \atbs_core_0.spike_memory_0.n2406_o[11]\ _00143_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[924]$_DFFE_PP0P_  clock_i _01874_ \atbs_core_0.spike_memory_0.n2406_o[12]\ _00146_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[925]$_DFFE_PP0P_  clock_i _01875_ \atbs_core_0.spike_memory_0.n2406_o[13]\ _00149_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[926]$_DFFE_PP0P_  clock_i _01876_ \atbs_core_0.spike_memory_0.n2406_o[14]\ _00007_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[927]$_DFFE_PP0P_  clock_i _01877_ \atbs_core_0.spike_memory_0.n2406_o[15]\ _00010_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[928]$_DFFE_PP0P_  clock_i _01878_ \atbs_core_0.spike_memory_0.n2406_o[16]\ _00013_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[929]$_DFFE_PP0P_  clock_i _01879_ \atbs_core_0.spike_memory_0.n2406_o[17]\ _00016_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[92]$_DFFE_PP0P_  clock_i _01880_ \atbs_core_0.spike_memory_0.n2362_o[16]\ _12858_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[930]$_DFFE_PP0P_  clock_i _01881_ \atbs_core_0.spike_memory_0.n2406_o[18]\ _00019_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[931]$_DFFE_PP0P_  clock_i _01882_ \atbs_core_0.spike_memory_0.n2407_o[0]\ _12857_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[932]$_DFFE_PP0P_  clock_i _01883_ \atbs_core_0.spike_memory_0.n2407_o[1]\ _12856_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[933]$_DFFE_PP0P_  clock_i _01884_ \atbs_core_0.spike_memory_0.n2407_o[2]\ _12855_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[934]$_DFFE_PP0P_  clock_i _01885_ \atbs_core_0.spike_memory_0.n2407_o[3]\ _12854_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[935]$_DFFE_PP0P_  clock_i _01886_ \atbs_core_0.spike_memory_0.n2407_o[4]\ _12853_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[936]$_DFFE_PP0P_  clock_i _01887_ \atbs_core_0.spike_memory_0.n2407_o[5]\ _12852_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[937]$_DFFE_PP0P_  clock_i _01888_ \atbs_core_0.spike_memory_0.n2407_o[6]\ _12851_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[938]$_DFFE_PP0P_  clock_i _01889_ \atbs_core_0.spike_memory_0.n2407_o[7]\ _12850_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[939]$_DFFE_PP0P_  clock_i _01890_ \atbs_core_0.spike_memory_0.n2407_o[8]\ _12849_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[93]$_DFFE_PP0P_  clock_i _01891_ \atbs_core_0.spike_memory_0.n2362_o[17]\ _12848_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[940]$_DFFE_PP0P_  clock_i _01892_ \atbs_core_0.spike_memory_0.n2407_o[9]\ _12847_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[941]$_DFFE_PP0P_  clock_i _01893_ \atbs_core_0.spike_memory_0.n2407_o[10]\ _12846_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[942]$_DFFE_PP0P_  clock_i _01894_ \atbs_core_0.spike_memory_0.n2407_o[11]\ _12845_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[943]$_DFFE_PP0P_  clock_i _01895_ \atbs_core_0.spike_memory_0.n2407_o[12]\ _12844_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[944]$_DFFE_PP0P_  clock_i _01896_ \atbs_core_0.spike_memory_0.n2407_o[13]\ _12843_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[945]$_DFFE_PP0P_  clock_i _01897_ \atbs_core_0.spike_memory_0.n2407_o[14]\ _12842_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[946]$_DFFE_PP0P_  clock_i _01898_ \atbs_core_0.spike_memory_0.n2407_o[15]\ _12841_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[947]$_DFFE_PP0P_  clock_i _01899_ \atbs_core_0.spike_memory_0.n2407_o[16]\ _12840_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[948]$_DFFE_PP0P_  clock_i _01900_ \atbs_core_0.spike_memory_0.n2407_o[17]\ _12839_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[949]$_DFFE_PP0P_  clock_i _01901_ \atbs_core_0.spike_memory_0.n2407_o[18]\ _12838_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[94]$_DFFE_PP0P_  clock_i _01902_ \atbs_core_0.spike_memory_0.n2362_o[18]\ _12837_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[950]$_DFFE_PP0P_  clock_i _01903_ \atbs_core_0.spike_memory_0.n2408_o[0]\ _12836_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[951]$_DFFE_PP0P_  clock_i _01904_ \atbs_core_0.spike_memory_0.n2408_o[1]\ _12835_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[952]$_DFFE_PP0P_  clock_i _01905_ \atbs_core_0.spike_memory_0.n2408_o[2]\ _12834_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[953]$_DFFE_PP0P_  clock_i _01906_ \atbs_core_0.spike_memory_0.n2408_o[3]\ _12833_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[954]$_DFFE_PP0P_  clock_i _01907_ \atbs_core_0.spike_memory_0.n2408_o[4]\ _12832_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[955]$_DFFE_PP0P_  clock_i _01908_ \atbs_core_0.spike_memory_0.n2408_o[5]\ _12831_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[956]$_DFFE_PP0P_  clock_i _01909_ \atbs_core_0.spike_memory_0.n2408_o[6]\ _12830_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[957]$_DFFE_PP0P_  clock_i _01910_ \atbs_core_0.spike_memory_0.n2408_o[7]\ _12829_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[958]$_DFFE_PP0P_  clock_i _01911_ \atbs_core_0.spike_memory_0.n2408_o[8]\ _12828_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[959]$_DFFE_PP0P_  clock_i _01912_ \atbs_core_0.spike_memory_0.n2408_o[9]\ _12827_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[95]$_DFFE_PP0P_  clock_i _01913_ \atbs_core_0.spike_memory_0.n2363_o[0]\ _12826_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[960]$_DFFE_PP0P_  clock_i _01914_ \atbs_core_0.spike_memory_0.n2408_o[10]\ _12825_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[961]$_DFFE_PP0P_  clock_i _01915_ \atbs_core_0.spike_memory_0.n2408_o[11]\ _12824_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[962]$_DFFE_PP0P_  clock_i _01916_ \atbs_core_0.spike_memory_0.n2408_o[12]\ _12823_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[963]$_DFFE_PP0P_  clock_i _01917_ \atbs_core_0.spike_memory_0.n2408_o[13]\ _12822_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[964]$_DFFE_PP0P_  clock_i _01918_ \atbs_core_0.spike_memory_0.n2408_o[14]\ _12821_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[965]$_DFFE_PP0P_  clock_i _01919_ \atbs_core_0.spike_memory_0.n2408_o[15]\ _12820_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[966]$_DFFE_PP0P_  clock_i _01920_ \atbs_core_0.spike_memory_0.n2408_o[16]\ _12819_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[967]$_DFFE_PP0P_  clock_i _01921_ \atbs_core_0.spike_memory_0.n2408_o[17]\ _12818_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[968]$_DFFE_PP0P_  clock_i _01922_ \atbs_core_0.spike_memory_0.n2408_o[18]\ _12817_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[969]$_DFFE_PP0P_  clock_i _01923_ \atbs_core_0.spike_memory_0.n2409_o[0]\ _12816_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[96]$_DFFE_PP0P_  clock_i _01924_ \atbs_core_0.spike_memory_0.n2363_o[1]\ _12815_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[970]$_DFFE_PP0P_  clock_i _01925_ \atbs_core_0.spike_memory_0.n2409_o[1]\ _12814_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[971]$_DFFE_PP0P_  clock_i _01926_ \atbs_core_0.spike_memory_0.n2409_o[2]\ _12813_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[972]$_DFFE_PP0P_  clock_i _01927_ \atbs_core_0.spike_memory_0.n2409_o[3]\ _12812_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[973]$_DFFE_PP0P_  clock_i _01928_ \atbs_core_0.spike_memory_0.n2409_o[4]\ _12811_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[974]$_DFFE_PP0P_  clock_i _01929_ \atbs_core_0.spike_memory_0.n2409_o[5]\ _12810_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[975]$_DFFE_PP0P_  clock_i _01930_ \atbs_core_0.spike_memory_0.n2409_o[6]\ _12809_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[976]$_DFFE_PP0P_  clock_i _01931_ \atbs_core_0.spike_memory_0.n2409_o[7]\ _12808_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[977]$_DFFE_PP0P_  clock_i _01932_ \atbs_core_0.spike_memory_0.n2409_o[8]\ _12807_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[978]$_DFFE_PP0P_  clock_i _01933_ \atbs_core_0.spike_memory_0.n2409_o[9]\ _12806_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[979]$_DFFE_PP0P_  clock_i _01934_ \atbs_core_0.spike_memory_0.n2409_o[10]\ _12805_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[97]$_DFFE_PP0P_  clock_i _01935_ \atbs_core_0.spike_memory_0.n2363_o[2]\ _12804_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[980]$_DFFE_PP0P_  clock_i _01936_ \atbs_core_0.spike_memory_0.n2409_o[11]\ _12803_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[981]$_DFFE_PP0P_  clock_i _01937_ \atbs_core_0.spike_memory_0.n2409_o[12]\ _12802_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[982]$_DFFE_PP0P_  clock_i _01938_ \atbs_core_0.spike_memory_0.n2409_o[13]\ _12801_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[983]$_DFFE_PP0P_  clock_i _01939_ \atbs_core_0.spike_memory_0.n2409_o[14]\ _12800_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[984]$_DFFE_PP0P_  clock_i _01940_ \atbs_core_0.spike_memory_0.n2409_o[15]\ _12799_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[985]$_DFFE_PP0P_  clock_i _01941_ \atbs_core_0.spike_memory_0.n2409_o[16]\ _12798_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[986]$_DFFE_PP0P_  clock_i _01942_ \atbs_core_0.spike_memory_0.n2409_o[17]\ _12797_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[987]$_DFFE_PP0P_  clock_i _01943_ \atbs_core_0.spike_memory_0.n2409_o[18]\ _12796_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[988]$_DFFE_PP0P_  clock_i _01944_ \atbs_core_0.spike_memory_0.n2410_o[0]\ _12795_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[989]$_DFFE_PP0P_  clock_i _01945_ \atbs_core_0.spike_memory_0.n2410_o[1]\ _12794_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[98]$_DFFE_PP0P_  clock_i _01946_ \atbs_core_0.spike_memory_0.n2363_o[3]\ _12793_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[990]$_DFFE_PP0P_  clock_i _01947_ \atbs_core_0.spike_memory_0.n2410_o[2]\ _12792_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[991]$_DFFE_PP0P_  clock_i _01948_ \atbs_core_0.spike_memory_0.n2410_o[3]\ _12791_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[992]$_DFFE_PP0P_  clock_i _01949_ \atbs_core_0.spike_memory_0.n2410_o[4]\ _12790_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[993]$_DFFE_PP0P_  clock_i _01950_ \atbs_core_0.spike_memory_0.n2410_o[5]\ _12789_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[994]$_DFFE_PP0P_  clock_i _01951_ \atbs_core_0.spike_memory_0.n2410_o[6]\ _12788_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[995]$_DFFE_PP0P_  clock_i _01952_ \atbs_core_0.spike_memory_0.n2410_o[7]\ _12787_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[996]$_DFFE_PP0P_  clock_i _01953_ \atbs_core_0.spike_memory_0.n2410_o[8]\ _12786_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[997]$_DFFE_PP0P_  clock_i _01954_ \atbs_core_0.spike_memory_0.n2410_o[9]\ _12785_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[998]$_DFFE_PP0P_  clock_i _01955_ \atbs_core_0.spike_memory_0.n2410_o[10]\ _12784_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[999]$_DFFE_PP0P_  clock_i _01956_ \atbs_core_0.spike_memory_0.n2410_o[11]\ _12783_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[99]$_DFFE_PP0P_  clock_i _01957_ \atbs_core_0.spike_memory_0.n2363_o[4]\ _12782_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2436_q[9]$_DFFE_PP0P_  clock_i _01958_ \atbs_core_0.spike_memory_0.n2358_o[9]\ _12781_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[0]$_DFFE_PP0P_  clock_i _01959_ \atbs_core_0.spike_memory_0.head[0]\ \atbs_core_0.spike_memory_0.n2306_o[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[1]$_DFFE_PP0P_  clock_i _01960_ \atbs_core_0.spike_memory_0.head[1]\ _12780_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[2]$_DFFE_PP0P_  clock_i _01961_ \atbs_core_0.spike_memory_0.head[2]\ _12779_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[3]$_DFFE_PP0P_  clock_i _01962_ \atbs_core_0.spike_memory_0.head[3]\ _12778_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[4]$_DFFE_PP0P_  clock_i _01963_ \atbs_core_0.spike_memory_0.head[4]\ _12777_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2437_q[5]$_DFFE_PP0P_  clock_i _01964_ \atbs_core_0.spike_memory_0.head[5]\ _12776_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[0]$_DFFE_PP0P_  clock_i _01965_ \atbs_core_0.spike_memory_0.n2438_q[0]\ \atbs_core_0.spike_memory_0.n2321_o[0]\ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[1]$_DFFE_PP0P_  clock_i _01966_ \atbs_core_0.spike_memory_0.n2438_q[1]\ _12775_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[2]$_DFFE_PP0P_  clock_i _01967_ \atbs_core_0.spike_memory_0.n2438_q[2]\ _12774_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[3]$_DFFE_PP0P_  clock_i _01968_ \atbs_core_0.spike_memory_0.n2438_q[3]\ _12773_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[4]$_DFFE_PP0P_  clock_i _01969_ \atbs_core_0.spike_memory_0.n2438_q[4]\ _12772_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2438_q[5]$_DFFE_PP0P_  clock_i _01970_ \atbs_core_0.spike_memory_0.n2438_q[5]\ _12771_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2439_q$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2304_o\ \atbs_core_0.spike_memory_0.n2439_q\ _12770_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[0]$_DFFE_PP0P_  clock_i _01971_ \atbs_core_0.spike_memory_0.a_data[0]\ _12769_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[10]$_DFFE_PP0P_  clock_i _01972_ \atbs_core_0.spike_memory_0.a_data[10]\ _12768_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[11]$_DFFE_PP0P_  clock_i _01973_ \atbs_core_0.spike_memory_0.a_data[11]\ _12767_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[12]$_DFFE_PP0P_  clock_i _01974_ \atbs_core_0.spike_memory_0.a_data[12]\ _12766_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[13]$_DFFE_PP0P_  clock_i _01975_ \atbs_core_0.spike_memory_0.a_data[13]\ _12765_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[14]$_DFFE_PP0P_  clock_i _01976_ \atbs_core_0.spike_memory_0.a_data[14]\ _12764_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[15]$_DFFE_PP0P_  clock_i _01977_ \atbs_core_0.spike_memory_0.a_data[15]\ _12763_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[16]$_DFFE_PP0P_  clock_i _01978_ \atbs_core_0.spike_memory_0.a_data[16]\ _12762_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[17]$_DFFE_PP0P_  clock_i _01979_ \atbs_core_0.spike_memory_0.a_data[17]\ _12761_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[18]$_DFFE_PP0P_  clock_i _01980_ \atbs_core_0.spike_memory_0.a_data[18]\ _12760_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[1]$_DFFE_PP0P_  clock_i _01981_ \atbs_core_0.spike_memory_0.a_data[1]\ _12759_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[2]$_DFFE_PP0P_  clock_i _01982_ \atbs_core_0.spike_memory_0.a_data[2]\ _12758_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[3]$_DFFE_PP0P_  clock_i _01983_ \atbs_core_0.spike_memory_0.a_data[3]\ _12757_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[4]$_DFFE_PP0P_  clock_i _01984_ \atbs_core_0.spike_memory_0.a_data[4]\ _12756_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[5]$_DFFE_PP0P_  clock_i _01985_ \atbs_core_0.spike_memory_0.a_data[5]\ _12755_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[6]$_DFFE_PP0P_  clock_i _01986_ \atbs_core_0.spike_memory_0.a_data[6]\ _12754_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[7]$_DFFE_PP0P_  clock_i _01987_ \atbs_core_0.spike_memory_0.a_data[7]\ _12753_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[8]$_DFFE_PP0P_  clock_i _01988_ \atbs_core_0.spike_memory_0.a_data[8]\ _12752_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2440_q[9]$_DFFE_PP0P_  clock_i _01989_ \atbs_core_0.spike_memory_0.a_data[9]\ _12751_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[0]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[0]\ \atbs_core_0.b_data[0]\ _12750_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[10]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[10]\ \atbs_core_0.b_data[10]\ _12749_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[11]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[11]\ \atbs_core_0.b_data[11]\ _12748_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[12]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[12]\ \atbs_core_0.b_data[12]\ _12747_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[13]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[13]\ \atbs_core_0.b_data[13]\ _12746_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[14]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[14]\ \atbs_core_0.b_data[14]\ _12745_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[15]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[15]\ \atbs_core_0.b_data[15]\ _12744_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[16]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[16]\ \atbs_core_0.b_data[16]\ _12743_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[17]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[17]\ \atbs_core_0.b_data[17]\ _12742_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[18]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[18]\ \atbs_core_0.b_data[18]\ _12741_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[1]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[1]\ \atbs_core_0.b_data[1]\ _12740_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[2]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[2]\ \atbs_core_0.b_data[2]\ _12739_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[3]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[3]\ \atbs_core_0.b_data[3]\ _12738_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[4]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[4]\ \atbs_core_0.b_data[4]\ _12737_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[5]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[5]\ \atbs_core_0.b_data[5]\ _12736_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[6]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[6]\ \atbs_core_0.b_data[6]\ _12735_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[7]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[7]\ \atbs_core_0.b_data[7]\ _12734_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[8]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[8]\ \atbs_core_0.b_data[8]\ _12733_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2441_q[9]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2550_o[9]\ \atbs_core_0.b_data[9]\ _12732_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2442_q[0]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2319_o\ \atbs_core_0.spike_memory_0.n2433_o\ _12731_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2442_q[1]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2433_o\ \atbs_core_0.spike_memory_0.n2431_o\ _12730_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2442_q[2]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2431_o\ \atbs_core_0.spike_memory_0.n2429_o\ _12729_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2442_q[3]$_DFF_PP0_  clock_i \atbs_core_0.spike_memory_0.n2429_o\ \atbs_core_0.memory2uart_0.read_strb_i\ _12728_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2444_q[0]$_DFFE_PP0P_  clock_i _01990_ \atbs_core_0.spike_memory_0.n2331_o\ _12727_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2444_q[1]$_DFFE_PP0P_  clock_i _01991_ \atbs_core_0.spike_memory_0.n2330_o\ _12726_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.spike_memory_0.n2444_q[2]$_DFFE_PP0P_  clock_i _01992_ \atbs_core_0.spike_memory_0.n2317_o\ _14572_ _00185_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_0.n1433_q[0]$_DFF_PN0_  clock_i _14577_ \atbs_core_0.sync_chain_0.n1426_o\ _14573_ reset_n_i VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_0.n1433_q[1]$_DFF_PN0_  clock_i \atbs_core_0.sync_chain_0.n1426_o\ \atbs_core_0.n66_o\ _12725_ reset_n_i VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1525_q[0]$_DFF_PP0_  clock_i comp_upper_i \atbs_core_0.sync_chain_1.buf[0]\ _12724_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1525_q[1]$_DFF_PP0_  clock_i comp_lower_i \atbs_core_0.sync_chain_1.buf[1]\ _12723_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1525_q[2]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_1.buf[0]\ \atbs_core_0.comp_upper_sync\ _12722_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_1.n1525_q[3]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_1.buf[1]\ \atbs_core_0.comp_lower_sync\ _12721_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_2.n1433_q[0]$_DFF_PP0_  clock_i trigger_start_sampling_i \atbs_core_0.sync_chain_2.n1426_o\ _12720_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.sync_chain_2.n1433_q[1]$_DFF_PP0_  clock_i \atbs_core_0.sync_chain_2.n1426_o\ \atbs_core_0.n72_o\ _12719_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[0]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[0]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[0]\ _00022_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[10]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[10]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[10]\ _00074_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[11]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[11]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[11]\ _00073_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[12]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[12]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[12]\ _00072_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[13]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[13]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[13]\ _00071_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[14]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[14]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[14]\ _00070_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[15]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[15]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[15]\ _00069_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[16]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[16]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[16]\ _00078_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[17]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[17]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[17]\ _00077_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[1]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[1]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[1]\ _00023_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[2]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[2]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[2]\ _00024_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[3]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[3]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[3]\ _00025_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[4]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[4]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[4]\ _00026_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[5]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[5]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[5]\ _00027_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[6]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[6]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[6]\ _00068_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[7]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[7]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[7]\ _00067_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[8]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[8]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[8]\ _00076_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2223_q[9]$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2218_o[9]\ \atbs_core_0.adaptive_ctrl_0.curr_time_i[9]\ _00075_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.time_measurement_0.n2224_q$_DFF_PP0_  clock_i \atbs_core_0.time_measurement_0.n2214_o\ \atbs_core_0.adaptive_ctrl_0.n1645_o\ _00100_ _00188_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3448_q[0]$_DFFE_PP0P_  clock_i _01993_ \atbs_core_0.uart_0.uart_rx_0.n3462_o\ _00063_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3448_q[1]$_DFFE_PP0P_  clock_i _01994_ \atbs_core_0.uart_0.uart_rx_0.n3456_o\ _12718_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3448_q[2]$_DFFE_PP0P_  clock_i _01995_ \atbs_core_0.uart_0.uart_rx_0.n3454_o\ _12717_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[0]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[0]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[0]\ _12716_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[1]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[1]\ _12715_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[2]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[2]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[2]\ _12714_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[3]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[3]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[3]\ _12713_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[4]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[4]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[4]\ _12712_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[5]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[5]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[5]\ _12711_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[6]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[6]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[6]\ _12710_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[7]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[7]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[7]\ _12709_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3449_q[8]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3401_o[8]\ \atbs_core_0.uart_0.uart_rx_0.baud_counter_value[8]\ _00057_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[0]$_DFFE_PP0P_  clock_i _01996_ \atbs_core_0.uart_0.uart_rx_0.n3472_o\ _12708_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[1]$_DFFE_PP0P_  clock_i _01997_ \atbs_core_0.uart_0.uart_rx_0.n3474_o\ _12707_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[2]$_DFFE_PP0P_  clock_i _01998_ \atbs_core_0.uart_0.uart_rx_0.n3476_o\ _12706_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[3]$_DFFE_PP0P_  clock_i _01999_ \atbs_core_0.uart_0.uart_rx_0.n3478_o\ _12705_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[4]$_DFFE_PP0P_  clock_i _02000_ \atbs_core_0.uart_0.uart_rx_0.n3480_o\ _12704_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[5]$_DFFE_PP0P_  clock_i _02001_ \atbs_core_0.uart_0.uart_rx_0.n3482_o\ _12703_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[6]$_DFFE_PP0P_  clock_i _02002_ \atbs_core_0.uart_0.uart_rx_0.n3484_o\ _12702_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3450_q[7]$_DFFE_PP0P_  clock_i _02003_ \atbs_core_0.uart_0.uart_rx_0.n3486_o\ _12701_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3451_q$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_rx_0.n3445_o\ \atbs_core_0.uart_0.rx_data_strb_o\ _12700_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3452_q[0]$_DFF_PP1_  clock_i _00189_ _14575_ \atbs_core_0.uart_0.uart_rx_0.n3399_o\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3452_q[1]$_DFF_PP0_  clock_i _00000_ \atbs_core_0.uart_0.uart_rx_0.n3384_o\ _12699_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3452_q[2]$_DFF_PP0_  clock_i _00001_ \atbs_core_0.uart_0.uart_rx_0.n3413_o\ _12698_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_rx_0.n3452_q[3]$_DFF_PP0_  clock_i _00002_ \atbs_core_0.uart_0.uart_rx_0.n3438_o\ _12697_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3344_q$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3341_o\ \atbs_core_0.memory2uart_0.tx_strb_i\ \atbs_core_0.spike_memory_0.n2333_o[0]\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3345_q[0]$_DFFE_PP0P_  clock_i _02004_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[0]\ _12696_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3345_q[1]$_DFFE_PP0P_  clock_i _02005_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[1]\ _12695_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3345_q[2]$_DFFE_PP0P_  clock_i _02006_ \atbs_core_0.uart_0.uart_tx_0.n3345_q[2]\ _00109_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[0]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[0]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[0]\ _12694_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[1]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[1]\ _12693_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[2]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[2]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[2]\ _12692_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[3]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[3]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[3]\ _12691_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[4]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[4]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[4]\ _12690_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[5]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[5]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[5]\ _12689_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[6]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[6]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[6]\ _12688_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[7]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[7]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[7]\ _12687_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3346_q[8]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3277_o[8]\ \atbs_core_0.uart_0.uart_tx_0.baud_counter_value[8]\ _12686_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3347_q[0]$_DFF_PP1_  clock_i _00190_ _14576_ \atbs_core_0.uart_0.uart_tx_0.n3286_o\ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3347_q[1]$_DFF_PP0_  clock_i \atbs_core_0.uart_0.uart_tx_0.n3331_o[2]\ \atbs_core_0.uart_0.uart_tx_0.n3323_o\ _00061_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3347_q[2]$_DFF_PP0_  clock_i _00003_ \atbs_core_0.uart_0.uart_tx_0.n3300_o\ _12685_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3347_q[3]$_DFF_PP0_  clock_i _00004_ \atbs_core_0.uart_0.uart_tx_0.n3295_o\ _12684_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1
X\atbs_core_0.uart_0.uart_tx_0.n3347_q[4]$_DFF_PP0_  clock_i _00005_ \atbs_core_0.uart_0.uart_tx_0.n3264_o\ _12683_ _00186_ VPWR 
+ VGND
+ sg13g2_dfrbp_1

.ends
.end
